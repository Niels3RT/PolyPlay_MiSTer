library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_char1 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_char1;

architecture rtl of rom_char1 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0000
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0008
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0010
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0018
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0020
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0028
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0030
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0038
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0040
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0048
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0050
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0058
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0060
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0068
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0070
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0078
         x"aa",  x"55",  x"aa",  x"55",  x"aa",  x"55",  x"aa",  x"55", -- 0080
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff", -- 0088
         x"3c",  x"24",  x"24",  x"66",  x"66",  x"66",  x"e7",  x"ff", -- 0090
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff", -- 0098
         x"42",  x"7e",  x"7e",  x"3c",  x"3c",  x"3c",  x"3c",  x"18", -- 00A0
         x"03",  x"1f",  x"ff",  x"c2",  x"c2",  x"ff",  x"1f",  x"03", -- 00A8
         x"ff",  x"ff",  x"ff",  x"18",  x"18",  x"ff",  x"ff",  x"ff", -- 00B0
         x"c0",  x"f8",  x"ff",  x"43",  x"43",  x"ff",  x"f8",  x"c0", -- 00B8
         x"1e",  x"0f",  x"07",  x"01",  x"07",  x"0f",  x"18",  x"00", -- 00C0
         x"46",  x"67",  x"ff",  x"ff",  x"9f",  x"33",  x"76",  x"cc", -- 00C8
         x"24",  x"3c",  x"bf",  x"ff",  x"ff",  x"ff",  x"dd",  x"c9", -- 00D0
         x"d0",  x"91",  x"bb",  x"ff",  x"ff",  x"ff",  x"b9",  x"88", -- 00D8
         x"f8",  x"f0",  x"c0",  x"30",  x"18",  x"c0",  x"e0",  x"70", -- 00E0
         x"08",  x"0c",  x"06",  x"0f",  x"3f",  x"07",  x"03",  x"01", -- 00E8
         x"95",  x"cd",  x"d7",  x"af",  x"ff",  x"ff",  x"ff",  x"ff", -- 00F0
         x"08",  x"70",  x"e0",  x"f0",  x"f8",  x"fc",  x"c0",  x"80", -- 00F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0100
         x"10",  x"10",  x"10",  x"10",  x"00",  x"10",  x"10",  x"00", -- 0108
         x"28",  x"28",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0110
         x"28",  x"7c",  x"28",  x"28",  x"7c",  x"28",  x"00",  x"00", -- 0118
         x"10",  x"3c",  x"50",  x"38",  x"14",  x"78",  x"10",  x"00", -- 0120
         x"52",  x"24",  x"08",  x"10",  x"24",  x"4a",  x"04",  x"00", -- 0128
         x"50",  x"50",  x"20",  x"52",  x"4a",  x"44",  x"3a",  x"00", -- 0130
         x"08",  x"10",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0138
         x"10",  x"20",  x"20",  x"20",  x"20",  x"10",  x"08",  x"00", -- 0140
         x"10",  x"08",  x"08",  x"08",  x"08",  x"10",  x"20",  x"00", -- 0148
         x"00",  x"44",  x"28",  x"7c",  x"28",  x"44",  x"00",  x"00", -- 0150
         x"00",  x"10",  x"10",  x"7c",  x"10",  x"10",  x"00",  x"00", -- 0158
         x"00",  x"00",  x"00",  x"00",  x"00",  x"18",  x"08",  x"10", -- 0160
         x"00",  x"00",  x"00",  x"7c",  x"00",  x"00",  x"00",  x"00", -- 0168
         x"00",  x"00",  x"00",  x"00",  x"00",  x"18",  x"18",  x"00", -- 0170
         x"02",  x"04",  x"08",  x"10",  x"20",  x"40",  x"80",  x"00", -- 0178
         x"18",  x"24",  x"42",  x"42",  x"42",  x"24",  x"18",  x"00", -- 0180
         x"10",  x"30",  x"10",  x"10",  x"10",  x"10",  x"38",  x"00", -- 0188
         x"38",  x"44",  x"04",  x"08",  x"10",  x"20",  x"7c",  x"00", -- 0190
         x"38",  x"44",  x"04",  x"18",  x"04",  x"44",  x"38",  x"00", -- 0198
         x"08",  x"10",  x"20",  x"48",  x"7c",  x"08",  x"08",  x"00", -- 01A0
         x"7c",  x"40",  x"40",  x"78",  x"04",  x"44",  x"38",  x"00", -- 01A8
         x"18",  x"20",  x"40",  x"78",  x"44",  x"44",  x"38",  x"00", -- 01B0
         x"7c",  x"04",  x"08",  x"10",  x"20",  x"20",  x"20",  x"00", -- 01B8
         x"38",  x"44",  x"44",  x"38",  x"44",  x"44",  x"38",  x"00", -- 01C0
         x"38",  x"44",  x"44",  x"3c",  x"04",  x"08",  x"30",  x"00", -- 01C8
         x"00",  x"00",  x"18",  x"18",  x"00",  x"18",  x"18",  x"00", -- 01D0
         x"00",  x"00",  x"18",  x"18",  x"00",  x"18",  x"08",  x"10", -- 01D8
         x"04",  x"08",  x"10",  x"20",  x"10",  x"08",  x"04",  x"00", -- 01E0
         x"00",  x"00",  x"7c",  x"00",  x"7c",  x"00",  x"00",  x"00", -- 01E8
         x"20",  x"10",  x"08",  x"04",  x"08",  x"10",  x"20",  x"00", -- 01F0
         x"44",  x"04",  x"08",  x"10",  x"10",  x"00",  x"10",  x"00", -- 01F8
         x"3c",  x"42",  x"4e",  x"52",  x"4c",  x"40",  x"3c",  x"00", -- 0200
         x"18",  x"24",  x"42",  x"7e",  x"42",  x"42",  x"42",  x"00", -- 0208
         x"78",  x"44",  x"44",  x"78",  x"44",  x"44",  x"78",  x"00", -- 0210
         x"1c",  x"22",  x"40",  x"40",  x"40",  x"22",  x"1c",  x"00", -- 0218
         x"78",  x"44",  x"42",  x"42",  x"42",  x"44",  x"78",  x"00", -- 0220
         x"7c",  x"40",  x"40",  x"78",  x"40",  x"40",  x"7c",  x"00", -- 0228
         x"7c",  x"40",  x"40",  x"78",  x"40",  x"40",  x"40",  x"00", -- 0230
         x"1c",  x"22",  x"40",  x"46",  x"42",  x"22",  x"1e",  x"00", -- 0238
         x"42",  x"42",  x"42",  x"7e",  x"42",  x"42",  x"42",  x"00", -- 0240
         x"38",  x"10",  x"10",  x"10",  x"10",  x"10",  x"38",  x"00", -- 0248
         x"1c",  x"08",  x"08",  x"08",  x"48",  x"48",  x"30",  x"00", -- 0250
         x"44",  x"48",  x"50",  x"60",  x"50",  x"48",  x"44",  x"00", -- 0258
         x"40",  x"40",  x"40",  x"40",  x"40",  x"40",  x"7c",  x"00", -- 0260
         x"82",  x"c6",  x"aa",  x"92",  x"92",  x"82",  x"82",  x"00", -- 0268
         x"42",  x"62",  x"52",  x"4a",  x"46",  x"42",  x"42",  x"00", -- 0270
         x"3c",  x"42",  x"42",  x"42",  x"42",  x"42",  x"3c",  x"00", -- 0278
         x"7c",  x"42",  x"42",  x"7c",  x"40",  x"40",  x"40",  x"00", -- 0280
         x"3c",  x"42",  x"42",  x"42",  x"4a",  x"44",  x"3a",  x"00", -- 0288
         x"7c",  x"42",  x"42",  x"7c",  x"48",  x"44",  x"42",  x"00", -- 0290
         x"3c",  x"42",  x"40",  x"3c",  x"02",  x"42",  x"3c",  x"00", -- 0298
         x"7c",  x"10",  x"10",  x"10",  x"10",  x"10",  x"10",  x"00", -- 02A0
         x"42",  x"42",  x"42",  x"42",  x"42",  x"42",  x"3c",  x"00", -- 02A8
         x"42",  x"42",  x"42",  x"42",  x"42",  x"24",  x"18",  x"00", -- 02B0
         x"82",  x"82",  x"92",  x"92",  x"92",  x"92",  x"6c",  x"00", -- 02B8
         x"82",  x"44",  x"28",  x"10",  x"28",  x"44",  x"82",  x"00", -- 02C0
         x"82",  x"44",  x"28",  x"10",  x"10",  x"10",  x"10",  x"00", -- 02C8
         x"7e",  x"04",  x"08",  x"10",  x"20",  x"40",  x"7e",  x"00", -- 02D0
         x"38",  x"20",  x"20",  x"20",  x"20",  x"20",  x"38",  x"00", -- 02D8
         x"80",  x"40",  x"20",  x"10",  x"08",  x"04",  x"02",  x"00", -- 02E0
         x"38",  x"08",  x"08",  x"08",  x"08",  x"08",  x"38",  x"00", -- 02E8
         x"10",  x"28",  x"44",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02F8
         x"62",  x"24",  x"28",  x"14",  x"2a",  x"44",  x"08",  x"0e", -- 0300
         x"00",  x"00",  x"34",  x"4c",  x"44",  x"4c",  x"34",  x"00", -- 0308
         x"40",  x"40",  x"58",  x"64",  x"44",  x"64",  x"58",  x"00", -- 0310
         x"00",  x"00",  x"38",  x"44",  x"40",  x"44",  x"38",  x"00", -- 0318
         x"04",  x"04",  x"34",  x"4c",  x"44",  x"4c",  x"34",  x"00", -- 0320
         x"00",  x"00",  x"38",  x"44",  x"78",  x"40",  x"3c",  x"00", -- 0328
         x"18",  x"24",  x"20",  x"70",  x"20",  x"20",  x"20",  x"00", -- 0330
         x"00",  x"00",  x"34",  x"4c",  x"44",  x"4c",  x"34",  x"04", -- 0338
         x"40",  x"40",  x"58",  x"64",  x"44",  x"44",  x"44",  x"00", -- 0340
         x"10",  x"00",  x"30",  x"10",  x"10",  x"10",  x"18",  x"00", -- 0348
         x"00",  x"08",  x"00",  x"18",  x"08",  x"08",  x"08",  x"48", -- 0350
         x"40",  x"40",  x"48",  x"50",  x"60",  x"50",  x"48",  x"00", -- 0358
         x"30",  x"10",  x"10",  x"10",  x"10",  x"14",  x"08",  x"00", -- 0360
         x"00",  x"00",  x"b6",  x"da",  x"92",  x"92",  x"92",  x"00", -- 0368
         x"00",  x"00",  x"58",  x"64",  x"44",  x"44",  x"44",  x"00", -- 0370
         x"00",  x"00",  x"38",  x"44",  x"44",  x"44",  x"38",  x"00", -- 0378
         x"00",  x"00",  x"58",  x"64",  x"44",  x"64",  x"58",  x"40", -- 0380
         x"00",  x"00",  x"34",  x"4c",  x"44",  x"4c",  x"34",  x"04", -- 0388
         x"00",  x"00",  x"58",  x"64",  x"40",  x"40",  x"40",  x"00", -- 0390
         x"00",  x"00",  x"3c",  x"40",  x"38",  x"04",  x"78",  x"00", -- 0398
         x"20",  x"20",  x"78",  x"20",  x"20",  x"24",  x"18",  x"00", -- 03A0
         x"00",  x"00",  x"44",  x"44",  x"44",  x"4c",  x"34",  x"00", -- 03A8
         x"00",  x"00",  x"44",  x"44",  x"44",  x"28",  x"10",  x"00", -- 03B0
         x"00",  x"00",  x"82",  x"92",  x"92",  x"92",  x"6c",  x"00", -- 03B8
         x"00",  x"00",  x"44",  x"28",  x"10",  x"28",  x"44",  x"00", -- 03C0
         x"00",  x"00",  x"44",  x"44",  x"44",  x"4c",  x"34",  x"04", -- 03C8
         x"00",  x"00",  x"7c",  x"08",  x"10",  x"20",  x"7c",  x"00", -- 03D0
         x"08",  x"10",  x"10",  x"20",  x"10",  x"10",  x"08",  x"00", -- 03D8
         x"10",  x"10",  x"10",  x"10",  x"10",  x"10",  x"10",  x"10", -- 03E0
         x"20",  x"10",  x"10",  x"08",  x"10",  x"10",  x"20",  x"00", -- 03E8
         x"18",  x"24",  x"20",  x"70",  x"20",  x"24",  x"7c",  x"00", -- 03F0
         x"24",  x"48",  x"12",  x"24",  x"48",  x"12",  x"24",  x"00"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
