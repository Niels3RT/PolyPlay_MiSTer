library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_7000 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_7000;

architecture rtl of rom1_7000 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"ff",  x"ff",  x"c3",  x"fb",  x"ff",  x"bf",  x"3e",  x"fc", -- 0000
         x"f0",  x"c0",  x"00",  x"00",  x"01",  x"07",  x"0f",  x"1f", -- 0008
         x"1f",  x"1f",  x"00",  x"00",  x"f2",  x"ff",  x"fe",  x"ff", -- 0010
         x"ff",  x"c1",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0018
         x"c0",  x"e0",  x"08",  x"00",  x"04",  x"1f",  x"07",  x"0f", -- 0020
         x"04",  x"00",  x"00",  x"00",  x"00",  x"c1",  x"c0",  x"f8", -- 0028
         x"fc",  x"7c",  x"3f",  x"0f",  x"03",  x"f0",  x"ff",  x"1f", -- 0030
         x"3f",  x"3f",  x"ff",  x"ff",  x"ff",  x"00",  x"80",  x"00", -- 0038
         x"80",  x"80",  x"80",  x"80",  x"00",  x"08",  x"00",  x"02", -- 0040
         x"07",  x"02",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0048
         x"fe",  x"fc",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0050
         x"08",  x"00",  x"02",  x"c3",  x"df",  x"ff",  x"fd",  x"7c", -- 0058
         x"3f",  x"0f",  x"03",  x"f1",  x"ff",  x"9f",  x"3f",  x"3f", -- 0060
         x"ff",  x"ff",  x"ff",  x"50",  x"00",  x"02",  x"00",  x"00", -- 0068
         x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"00",  x"f0", -- 0070
         x"f0",  x"0f",  x"0f",  x"00",  x"00",  x"00",  x"10",  x"00", -- 0078
         x"02",  x"18",  x"3c",  x"7e",  x"ff",  x"7e",  x"3c",  x"18", -- 0080
         x"00",  x"18",  x"3c",  x"7e",  x"ff",  x"7e",  x"3c",  x"18", -- 0088
         x"00",  x"20",  x"00",  x"03",  x"00",  x"03",  x"00",  x"00", -- 0090
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0098
         x"06",  x"3f",  x"3f",  x"06",  x"00",  x"0c",  x"00",  x"00", -- 00A0
         x"00",  x"c0",  x"c0",  x"00",  x"08",  x"00",  x"01",  x"00", -- 00A8
         x"00",  x"03",  x"00",  x"00",  x"00",  x"00",  x"00",  x"08", -- 00B0
         x"00",  x"01",  x"00",  x"00",  x"0c",  x"00",  x"00",  x"00", -- 00B8
         x"00",  x"00",  x"08",  x"00",  x"02",  x"00",  x"00",  x"00", -- 00C0
         x"00",  x"06",  x"3f",  x"3f",  x"06",  x"00",  x"0c",  x"00", -- 00C8
         x"00",  x"00",  x"c0",  x"c0",  x"00",  x"20",  x"00",  x"03", -- 00D0
         x"01",  x"01",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00D8
         x"00",  x"00",  x"00",  x"06",  x"06",  x"1f",  x"1f",  x"06", -- 00E0
         x"08",  x"08",  x"00",  x"00",  x"00",  x"80",  x"80",  x"00", -- 00E8
         x"08",  x"00",  x"03",  x"00",  x"00",  x"01",  x"01",  x"00", -- 00F0
         x"00",  x"00",  x"00",  x"06",  x"00",  x"00",  x"00",  x"00", -- 00F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"08",  x"08",  x"00", -- 0100
         x"00",  x"00",  x"00",  x"08",  x"00",  x"02",  x"00",  x"00", -- 0108
         x"00",  x"06",  x"06",  x"1f",  x"1f",  x"06",  x"08",  x"08", -- 0110
         x"00",  x"00",  x"00",  x"80",  x"80",  x"00",  x"08",  x"00", -- 0118
         x"01",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"04", -- 0120
         x"0c",  x"10",  x"00",  x"03",  x"00",  x"00",  x"00",  x"00", -- 0128
         x"00",  x"18",  x"08",  x"00",  x"00",  x"00",  x"00",  x"10", -- 0130
         x"3c",  x"1f",  x"1f",  x"0b",  x"00",  x"00",  x"00",  x"00", -- 0138
         x"00",  x"80",  x"03",  x"82",  x"10",  x"00",  x"01",  x"00", -- 0140
         x"00",  x"00",  x"00",  x"06",  x"04",  x"00",  x"00",  x"10", -- 0148
         x"00",  x"02",  x"00",  x"00",  x"00",  x"10",  x"3c",  x"1f", -- 0150
         x"1f",  x"0b",  x"00",  x"00",  x"00",  x"00",  x"00",  x"80", -- 0158
         x"03",  x"82",  x"10",  x"00",  x"01",  x"00",  x"00",  x"00", -- 0160
         x"00",  x"00",  x"00",  x"20",  x"30",  x"10",  x"00",  x"03", -- 0168
         x"00",  x"00",  x"00",  x"00",  x"00",  x"01",  x"c0",  x"41", -- 0170
         x"00",  x"00",  x"00",  x"08",  x"3c",  x"f8",  x"f8",  x"d0", -- 0178
         x"00",  x"00",  x"00",  x"00",  x"00",  x"18",  x"10",  x"00", -- 0180
         x"10",  x"00",  x"01",  x"00",  x"00",  x"00",  x"00",  x"60", -- 0188
         x"20",  x"00",  x"00",  x"08",  x"00",  x"03",  x"00",  x"00", -- 0190
         x"00",  x"00",  x"00",  x"01",  x"c0",  x"41",  x"00",  x"00", -- 0198
         x"00",  x"08",  x"3c",  x"f8",  x"f8",  x"d0",  x"00",  x"00", -- 01A0
         x"00",  x"00",  x"00",  x"03",  x"00",  x"00",  x"08",  x"00", -- 01A8
         x"01",  x"00",  x"00",  x"00",  x"00",  x"00",  x"0c",  x"00", -- 01B0
         x"00",  x"08",  x"00",  x"03",  x"00",  x"00",  x"00",  x"00", -- 01B8
         x"00",  x"00",  x"03",  x"00",  x"06",  x"3f",  x"3f",  x"06", -- 01C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"c0",  x"c0",  x"00", -- 01C8
         x"00",  x"00",  x"0c",  x"00",  x"28",  x"00",  x"02",  x"06", -- 01D0
         x"3f",  x"3f",  x"06",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01D8
         x"c0",  x"c0",  x"00",  x"00",  x"00",  x"0c",  x"00",  x"28", -- 01E0
         x"00",  x"03",  x"10",  x"10",  x"00",  x"00",  x"00",  x"01", -- 01E8
         x"01",  x"00",  x"00",  x"00",  x"00",  x"60",  x"60",  x"f8", -- 01F0
         x"f8",  x"60",  x"80",  x"80",  x"00",  x"00",  x"00",  x"00", -- 01F8
         x"00",  x"00",  x"08",  x"00",  x"05",  x"00",  x"00",  x"10", -- 0200
         x"10",  x"00",  x"00",  x"00",  x"00",  x"60",  x"00",  x"00", -- 0208
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"80", -- 0210
         x"80",  x"00",  x"00",  x"00",  x"00",  x"10",  x"10",  x"00", -- 0218
         x"00",  x"00",  x"01",  x"01",  x"00",  x"00",  x"00",  x"00", -- 0220
         x"60",  x"60",  x"f8",  x"f8",  x"60",  x"08",  x"00",  x"02", -- 0228
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"01", -- 0230
         x"00",  x"00",  x"40",  x"c0",  x"00",  x"00",  x"00",  x"00", -- 0238
         x"08",  x"00",  x"04",  x"00",  x"01",  x"00",  x"00",  x"00", -- 0240
         x"00",  x"00",  x"00",  x"03",  x"81",  x"81",  x"00",  x"00", -- 0248
         x"00",  x"00",  x"00",  x"c0",  x"f8",  x"f0",  x"b8",  x"00", -- 0250
         x"00",  x"00",  x"00",  x"00",  x"00",  x"30",  x"20",  x"00", -- 0258
         x"00",  x"00",  x"00",  x"10",  x"00",  x"01",  x"60",  x"40", -- 0260
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"08",  x"00", -- 0268
         x"02",  x"03",  x"81",  x"81",  x"00",  x"00",  x"00",  x"00", -- 0270
         x"00",  x"c0",  x"f8",  x"f0",  x"b8",  x"00",  x"00",  x"00", -- 0278
         x"00",  x"08",  x"00",  x"02",  x"00",  x"00",  x"02",  x"03", -- 0280
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0288
         x"00",  x"00",  x"00",  x"80",  x"08",  x"00",  x"04",  x"00", -- 0290
         x"00",  x"0c",  x"04",  x"00",  x"00",  x"00",  x"00",  x"03", -- 0298
         x"1f",  x"0f",  x"1d",  x"00",  x"00",  x"00",  x"00",  x"c0", -- 02A0
         x"81",  x"81",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02A8
         x"80",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"08", -- 02B0
         x"00",  x"01",  x"06",  x"02",  x"00",  x"00",  x"00",  x"00", -- 02B8
         x"00",  x"00",  x"10",  x"00",  x"02",  x"03",  x"1f",  x"0f", -- 02C0
         x"1d",  x"00",  x"00",  x"00",  x"00",  x"c0",  x"81",  x"81", -- 02C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"58",  x"00",  x"02", -- 02D0
         x"00",  x"f0",  x"f0",  x"0f",  x"0f",  x"00",  x"00",  x"00", -- 02D8
         x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02E0
         x"10",  x"00",  x"01",  x"18",  x"3c",  x"7e",  x"ff",  x"7e", -- 02E8
         x"3c",  x"18",  x"00",  x"3e",  x"ff",  x"ff",  x"ff",  x"ff", -- 02F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02F8
         x"00",  x"00",  x"03",  x"00",  x"00",  x"00",  x"3f",  x"7f", -- 0300
         x"ff",  x"ff",  x"ff",  x"f9",  x"e0",  x"00",  x"c0",  x"f0", -- 0308
         x"f0",  x"f0",  x"fc",  x"f0",  x"70",  x"08",  x"00",  x"03", -- 0310
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"03",  x"00", -- 0318
         x"e0",  x"f0",  x"f0",  x"e0",  x"e0",  x"f9",  x"ff",  x"ff", -- 0320
         x"70",  x"f0",  x"f0",  x"70",  x"70",  x"f0",  x"fc",  x"f0", -- 0328
         x"10",  x"00",  x"02",  x"ff",  x"7f",  x"3f",  x"00",  x"00", -- 0330
         x"00",  x"00",  x"00",  x"f0",  x"e0",  x"c0",  x"00",  x"00", -- 0338
         x"00",  x"00",  x"00",  x"08",  x"00",  x"02",  x"e6",  x"ff", -- 0340
         x"ff",  x"e6",  x"e0",  x"f9",  x"ff",  x"ff",  x"70",  x"f0", -- 0348
         x"f0",  x"70",  x"70",  x"f0",  x"fc",  x"f0",  x"20",  x"00", -- 0350
         x"0a",  x"00",  x"00",  x"01",  x"03",  x"07",  x"07",  x"07", -- 0358
         x"07",  x"10",  x"10",  x"ff",  x"ff",  x"fc",  x"f0",  x"f0", -- 0360
         x"fc",  x"00",  x"00",  x"ff",  x"ff",  x"63",  x"00",  x"00", -- 0368
         x"63",  x"80",  x"80",  x"f8",  x"fc",  x"fe",  x"fe",  x"fe", -- 0370
         x"fe",  x"03",  x"01",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0378
         x"00",  x"ff",  x"ff",  x"10",  x"10",  x"00",  x"00",  x"00", -- 0380
         x"00",  x"ff",  x"ff",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0388
         x"00",  x"fc",  x"f8",  x"80",  x"80",  x"00",  x"00",  x"00", -- 0390
         x"00",  x"10",  x"10",  x"ff",  x"ff",  x"fc",  x"f1",  x"f1", -- 0398
         x"fc",  x"00",  x"00",  x"ff",  x"ff",  x"63",  x"f8",  x"f8", -- 03A0
         x"63",  x"08",  x"00",  x"07",  x"00",  x"00",  x"00",  x"00", -- 03A8
         x"00",  x"00",  x"03",  x"07",  x"00",  x"00",  x"4f",  x"ff", -- 03B0
         x"7f",  x"ff",  x"ff",  x"83",  x"00",  x"00",  x"80",  x"e0", -- 03B8
         x"f0",  x"f8",  x"f8",  x"f8",  x"00",  x"01",  x"00",  x"01", -- 03C0
         x"01",  x"01",  x"01",  x"00",  x"0f",  x"ff",  x"f8",  x"fc", -- 03C8
         x"fc",  x"ff",  x"ff",  x"ff",  x"83",  x"03",  x"1f",  x"3f", -- 03D0
         x"3e",  x"fc",  x"f0",  x"c0",  x"f8",  x"e0",  x"f0",  x"20", -- 03D8
         x"00",  x"00",  x"00",  x"00",  x"08",  x"00",  x"02",  x"7f", -- 03E0
         x"3f",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"e0", -- 03E8
         x"40",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"08", -- 03F0
         x"00",  x"05",  x"0f",  x"ff",  x"f9",  x"fc",  x"fc",  x"ff"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
