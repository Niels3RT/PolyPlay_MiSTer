library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_5c00 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_5c00;

architecture rtl of rom1_5c00 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"e4",  x"20",  x"20",  x"ca",  x"cc",  x"e0",  x"e2",  x"e4", -- 0000
         x"20",  x"f6",  x"f8",  x"ca",  x"fa",  x"e0",  x"e2",  x"e4", -- 0008
         x"20",  x"40",  x"00",  x"40",  x"18",  x"41",  x"20",  x"c1", -- 0010
         x"18",  x"00",  x"00",  x"40",  x"08",  x"3f",  x"10",  x"bf", -- 0018
         x"08",  x"00",  x"00",  x"40",  x"18",  x"41",  x"20",  x"c1", -- 0020
         x"18",  x"00",  x"00",  x"40",  x"08",  x"3f",  x"10",  x"bf", -- 0028
         x"08",  x"00",  x"00",  x"00",  x"00",  x"00",  x"80",  x"00", -- 0030
         x"ff",  x"a7",  x"a1",  x"a9",  x"a3",  x"ab",  x"a5",  x"20", -- 0038
         x"20",  x"00",  x"02",  x"ff",  x"03",  x"80",  x"00",  x"90", -- 0040
         x"94",  x"02",  x"09",  x"01",  x"38",  x"01",  x"18",  x"00", -- 0048
         x"0c",  x"83",  x"87",  x"01",  x"0c",  x"83",  x"87",  x"01", -- 0050
         x"0c",  x"83",  x"87",  x"01",  x"30",  x"c4",  x"00",  x"08", -- 0058
         x"83",  x"87",  x"01",  x"18",  x"93",  x"00",  x"01",  x"20", -- 0060
         x"04",  x"28",  x"01",  x"20",  x"04",  x"28",  x"00",  x"00", -- 0068
         x"00",  x"05",  x"03",  x"0f",  x"3f",  x"7f",  x"7f",  x"ff", -- 0070
         x"ff",  x"ff",  x"c0",  x"f0",  x"fc",  x"fe",  x"fe",  x"ff", -- 0078
         x"ff",  x"ff",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0080
         x"00",  x"00",  x"ff",  x"7f",  x"7f",  x"3f",  x"0f",  x"03", -- 0088
         x"07",  x"00",  x"ff",  x"fe",  x"fe",  x"fc",  x"f0",  x"c0", -- 0090
         x"e0",  x"00",  x"30",  x"02",  x"06",  x"ff",  x"ff",  x"ff", -- 0098
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"00",  x"00", -- 00A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff", -- 00B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"00",  x"00", -- 00B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff", -- 00C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"20",  x"01",  x"01", -- 00C8
         x"00",  x"00",  x"00",  x"03",  x"0e",  x"00",  x"00",  x"00", -- 00D0
         x"70",  x"00",  x"05",  x"01",  x"03",  x"07",  x"07",  x"03", -- 00D8
         x"01",  x"07",  x"3f",  x"e0",  x"f8",  x"9c",  x"fc",  x"f8", -- 00E0
         x"e0",  x"f1",  x"fd",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00E8
         x"00",  x"00",  x"00",  x"7f",  x"71",  x"78",  x"3e",  x"0f", -- 00F0
         x"03",  x"00",  x"00",  x"ff",  x"ff",  x"07",  x"1e",  x"fc", -- 00F8
         x"e0",  x"00",  x"00",  x"30",  x"00",  x"05",  x"07",  x"1f", -- 0100
         x"39",  x"3f",  x"1f",  x"07",  x"8f",  x"bf",  x"80",  x"c0", -- 0108
         x"e0",  x"e0",  x"c0",  x"80",  x"e0",  x"fc",  x"00",  x"00", -- 0110
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff", -- 0118
         x"e0",  x"78",  x"3f",  x"07",  x"00",  x"00",  x"fe",  x"8e", -- 0120
         x"1e",  x"7c",  x"f0",  x"c0",  x"00",  x"00",  x"30",  x"00", -- 0128
         x"05",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"03", -- 0130
         x"07",  x"00",  x"00",  x"00",  x"00",  x"00",  x"80",  x"e0", -- 0138
         x"f0",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0140
         x"00",  x"07",  x"03",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0148
         x"00",  x"f0",  x"e0",  x"80",  x"00",  x"00",  x"00",  x"00", -- 0150
         x"00",  x"30",  x"00",  x"1f",  x"60",  x"60",  x"60",  x"60", -- 0158
         x"60",  x"60",  x"60",  x"60",  x"00",  x"00",  x"00",  x"03", -- 0160
         x"07",  x"1f",  x"ff",  x"ff",  x"00",  x"00",  x"80",  x"80", -- 0168
         x"80",  x"80",  x"90",  x"90",  x"00",  x"55",  x"aa",  x"55", -- 0170
         x"aa",  x"55",  x"aa",  x"55",  x"00",  x"00",  x"00",  x"00", -- 0178
         x"00",  x"00",  x"00",  x"00",  x"00",  x"07",  x"1f",  x"3c", -- 0180
         x"3c",  x"3f",  x"1f",  x"0f",  x"00",  x"00",  x"e0",  x"f0", -- 0188
         x"f0",  x"f0",  x"e0",  x"80",  x"00",  x"00",  x"00",  x"ff", -- 0190
         x"ff",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0198
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"18",  x"18", -- 01A0
         x"18",  x"18",  x"18",  x"7e",  x"18",  x"18",  x"18",  x"ff", -- 01A8
         x"ff",  x"18",  x"18",  x"18",  x"ff",  x"ff",  x"ff",  x"ff", -- 01B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 01B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"00",  x"00",  x"00", -- 01C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"07",  x"0f", -- 01C8
         x"0f",  x"0f",  x"07",  x"01",  x"00",  x"e0",  x"f8",  x"3c", -- 01D0
         x"3c",  x"fc",  x"f8",  x"f0",  x"fc",  x"fe",  x"ff",  x"7f", -- 01D8
         x"3f",  x"0f",  x"03",  x"00",  x"7e",  x"ff",  x"7e",  x"7e", -- 01E0
         x"ff",  x"ff",  x"ff",  x"00",  x"3f",  x"7f",  x"ff",  x"fe", -- 01E8
         x"fc",  x"f0",  x"c0",  x"00",  x"00",  x"00",  x"70",  x"f0", -- 01F0
         x"b8",  x"3e",  x"1f",  x"0f",  x"7e",  x"99",  x"ff",  x"81", -- 01F8
         x"42",  x"e7",  x"ff",  x"ff",  x"00",  x"00",  x"0e",  x"0f", -- 0200
         x"1d",  x"7c",  x"f8",  x"f0",  x"07",  x"03",  x"01",  x"01", -- 0208
         x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff",  x"ff", -- 0210
         x"bd",  x"18",  x"00",  x"00",  x"e0",  x"c0",  x"80",  x"80", -- 0218
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0220
         x"03",  x"07",  x"17",  x"7f",  x"0f",  x"1f",  x"7f",  x"fe", -- 0228
         x"fe",  x"fc",  x"f8",  x"f0",  x"f0",  x"f8",  x"fe",  x"7f", -- 0230
         x"7f",  x"3f",  x"1f",  x"0f",  x"00",  x"00",  x"00",  x"00", -- 0238
         x"c0",  x"e0",  x"f8",  x"fc",  x"00",  x"00",  x"c0",  x"e0", -- 0240
         x"e0",  x"e0",  x"c0",  x"80",  x"00",  x"00",  x"03",  x"07", -- 0248
         x"07",  x"07",  x"03",  x"01",  x"30",  x"00",  x"03",  x"00", -- 0250
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0258
         x"00",  x"00",  x"00",  x"00",  x"00",  x"03",  x"00",  x"00", -- 0260
         x"00",  x"00",  x"00",  x"00",  x"00",  x"c0",  x"00",  x"30", -- 0268
         x"00",  x"05",  x"81",  x"63",  x"1f",  x"37",  x"c3",  x"01", -- 0270
         x"07",  x"3f",  x"e0",  x"f8",  x"9c",  x"fc",  x"f8",  x"e0", -- 0278
         x"f1",  x"fd",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0280
         x"00",  x"00",  x"7f",  x"71",  x"78",  x"3e",  x"0f",  x"03", -- 0288
         x"00",  x"0f",  x"ff",  x"ff",  x"07",  x"1e",  x"fc",  x"f8", -- 0290
         x"18",  x"f8",  x"30",  x"00",  x"05",  x"07",  x"1f",  x"39", -- 0298
         x"3f",  x"1f",  x"07",  x"8f",  x"bf",  x"81",  x"c6",  x"f8", -- 02A0
         x"ec",  x"c3",  x"80",  x"e0",  x"fc",  x"00",  x"00",  x"00", -- 02A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"e0", -- 02B0
         x"78",  x"3f",  x"1f",  x"18",  x"1f",  x"fe",  x"8e",  x"1e", -- 02B8
         x"7c",  x"f0",  x"c0",  x"00",  x"f0",  x"30",  x"00",  x"05", -- 02C0
         x"00",  x"00",  x"00",  x"39",  x"3d",  x"1f",  x"0f",  x"7f", -- 02C8
         x"00",  x"00",  x"80",  x"ce",  x"de",  x"fc",  x"f8",  x"ff", -- 02D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02D8
         x"ff",  x"0f",  x"1f",  x"3d",  x"39",  x"00",  x"00",  x"00", -- 02E0
         x"ff",  x"f8",  x"fc",  x"de",  x"ce",  x"80",  x"00",  x"00", -- 02E8
         x"50",  x"00",  x"1d",  x"60",  x"60",  x"60",  x"60",  x"60", -- 02F0
         x"60",  x"60",  x"60",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0300
         x"00",  x"00",  x"00",  x"00",  x"07",  x"1f",  x"3c",  x"3c", -- 0308
         x"3f",  x"1f",  x"0f",  x"00",  x"01",  x"e3",  x"f6",  x"fc", -- 0310
         x"fc",  x"e6",  x"83",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0318
         x"00",  x"00",  x"00",  x"00",  x"18",  x"3c",  x"7e",  x"7e", -- 0320
         x"3c",  x"18",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0328
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0330
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0338
         x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0340
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0348
         x"ff",  x"ff",  x"ff",  x"00",  x"80",  x"c7",  x"6f",  x"3f", -- 0350
         x"3f",  x"67",  x"c1",  x"00",  x"e0",  x"f8",  x"3c",  x"3c", -- 0358
         x"fc",  x"f8",  x"f0",  x"fc",  x"fe",  x"ff",  x"7f",  x"3f", -- 0360
         x"0f",  x"03",  x"00",  x"7e",  x"ff",  x"7e",  x"7e",  x"ff", -- 0368
         x"ff",  x"ff",  x"7e",  x"3f",  x"7f",  x"ff",  x"fe",  x"fc", -- 0370
         x"f0",  x"c0",  x"00",  x"00",  x"00",  x"70",  x"f0",  x"b8", -- 0378
         x"3e",  x"1f",  x"0f",  x"7e",  x"99",  x"ff",  x"ff",  x"7e", -- 0380
         x"ff",  x"ff",  x"ff",  x"00",  x"00",  x"0e",  x"0f",  x"1d", -- 0388
         x"7c",  x"f8",  x"f0",  x"07",  x"03",  x"01",  x"01",  x"00", -- 0390
         x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0398
         x"5a",  x"42",  x"e7",  x"e0",  x"c0",  x"80",  x"80",  x"00", -- 03A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"03", -- 03A8
         x"07",  x"17",  x"7f",  x"0f",  x"1f",  x"7f",  x"fe",  x"fe", -- 03B0
         x"fc",  x"f8",  x"f0",  x"f0",  x"f8",  x"fe",  x"7f",  x"7f", -- 03B8
         x"3f",  x"1f",  x"0f",  x"00",  x"00",  x"00",  x"00",  x"c0", -- 03C0
         x"e0",  x"f8",  x"fc",  x"00",  x"00",  x"c0",  x"e0",  x"ff", -- 03C8
         x"ff",  x"c0",  x"80",  x"00",  x"00",  x"03",  x"07",  x"ff", -- 03D0
         x"ff",  x"03",  x"01",  x"0c",  x"ff",  x"ff",  x"ff",  x"ff", -- 03D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
