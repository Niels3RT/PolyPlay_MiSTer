library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_8c00 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_8c00;

architecture rtl of rom1_8c00 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"20", -- 0000
         x"50",  x"55",  x"4e",  x"4b",  x"54",  x"45",  x"3a",  x"20", -- 0008
         x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"20", -- 0010
         x"53",  x"50",  x"49",  x"45",  x"4c",  x"3a",  x"20",  x"3d", -- 0018
         x"3d",  x"3d",  x"3d",  x"25",  x"20",  x"57",  x"41",  x"53", -- 0020
         x"53",  x"45",  x"52",  x"53",  x"54",  x"26",  x"3a",  x"20", -- 0028
         x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"57",  x"20",  x"41", -- 0030
         x"20",  x"53",  x"20",  x"53",  x"20",  x"45",  x"20",  x"52", -- 0038
         x"20",  x"52",  x"20",  x"4f",  x"20",  x"48",  x"20",  x"52", -- 0040
         x"20",  x"42",  x"20",  x"52",  x"20",  x"55",  x"20",  x"43", -- 0048
         x"20",  x"48",  x"49",  x"4d",  x"20",  x"4f",  x"42",  x"45", -- 0050
         x"52",  x"45",  x"4e",  x"20",  x"5a",  x"49",  x"4d",  x"4d", -- 0058
         x"45",  x"52",  x"20",  x"49",  x"53",  x"54",  x"20",  x"45", -- 0060
         x"49",  x"4e",  x"20",  x"57",  x"41",  x"53",  x"53",  x"45", -- 0068
         x"52",  x"52",  x"4f",  x"48",  x"52",  x"20",  x"47",  x"45", -- 0070
         x"2d",  x"00",  x"00",  x"00",  x"00",  x"00",  x"50",  x"4c", -- 0078
         x"41",  x"54",  x"5a",  x"54",  x"2e",  x"20",  x"44",  x"55", -- 0080
         x"52",  x"43",  x"48",  x"20",  x"44",  x"41",  x"53",  x"20", -- 0088
         x"41",  x"55",  x"46",  x"46",  x"41",  x"4e",  x"47",  x"45", -- 0090
         x"4e",  x"20",  x"44",  x"45",  x"52",  x"20",  x"54",  x"52", -- 0098
         x"4f",  x"50",  x"46",  x"45",  x"4e",  x"20",  x"4d",  x"49", -- 00A0
         x"54",  x"00",  x"44",  x"45",  x"4d",  x"20",  x"45",  x"49", -- 00A8
         x"4d",  x"45",  x"52",  x"20",  x"4b",  x"41",  x"4e",  x"4e", -- 00B0
         x"20",  x"4d",  x"41",  x"4e",  x"20",  x"56",  x"45",  x"52", -- 00B8
         x"48",  x"49",  x"4e",  x"44",  x"45",  x"52",  x"4e",  x"2c", -- 00C0
         x"20",  x"44",  x"41",  x"53",  x"53",  x"20",  x"44",  x"45", -- 00C8
         x"52",  x"20",  x"57",  x"41",  x"53",  x"2d",  x"53",  x"45", -- 00D0
         x"52",  x"53",  x"54",  x"41",  x"4e",  x"44",  x"20",  x"53", -- 00D8
         x"54",  x"45",  x"49",  x"47",  x"54",  x"2e",  x"20",  x"44", -- 00E0
         x"45",  x"4e",  x"20",  x"45",  x"49",  x"4d",  x"45",  x"52", -- 00E8
         x"20",  x"4b",  x"41",  x"4e",  x"4e",  x"20",  x"4d",  x"41", -- 00F0
         x"4e",  x"20",  x"5a",  x"55",  x"4d",  x"00",  x"00",  x"00", -- 00F8
         x"00",  x"00",  x"4b",  x"45",  x"4c",  x"4c",  x"45",  x"52", -- 0100
         x"46",  x"45",  x"4e",  x"53",  x"54",  x"45",  x"52",  x"20", -- 0108
         x"41",  x"55",  x"53",  x"53",  x"43",  x"48",  x"55",  x"45", -- 0110
         x"54",  x"54",  x"45",  x"4e",  x"20",  x"28",  x"53",  x"50", -- 0118
         x"49",  x"45",  x"4c",  x"4b",  x"4e",  x"4f",  x"50",  x"46", -- 0120
         x"29",  x"2e",  x"00",  x"00",  x"00",  x"00",  x"49",  x"53", -- 0128
         x"54",  x"20",  x"44",  x"45",  x"52",  x"20",  x"45",  x"49", -- 0130
         x"4d",  x"45",  x"52",  x"20",  x"56",  x"4f",  x"4c",  x"4c", -- 0138
         x"20",  x"42",  x"45",  x"4b",  x"4f",  x"4d",  x"4d",  x"54", -- 0140
         x"20",  x"4d",  x"41",  x"4e",  x"20",  x"4b",  x"45",  x"49", -- 0148
         x"4e",  x"45",  x"20",  x"50",  x"55",  x"4e",  x"4b",  x"54", -- 0150
         x"45",  x"2e",  x"50",  x"55",  x"4e",  x"4b",  x"54",  x"45", -- 0158
         x"57",  x"45",  x"52",  x"54",  x"55",  x"4e",  x"47",  x"3a", -- 0160
         x"57",  x"41",  x"53",  x"53",  x"45",  x"52",  x"53",  x"54", -- 0168
         x"41",  x"4e",  x"44",  x"20",  x"5a",  x"55",  x"20",  x"48", -- 0170
         x"4f",  x"43",  x"48",  x"3a",  x"20",  x"20",  x"20",  x"20", -- 0178
         x"20",  x"20",  x"20",  x"2d",  x"31",  x"20",  x"53",  x"50", -- 0180
         x"49",  x"45",  x"4c",  x"41",  x"55",  x"46",  x"47",  x"45", -- 0188
         x"46",  x"41",  x"4e",  x"47",  x"45",  x"4e",  x"45",  x"52", -- 0190
         x"20",  x"54",  x"52",  x"4f",  x"50",  x"46",  x"45",  x"4e", -- 0198
         x"3a",  x"20",  x"20",  x"20",  x"20",  x"20",  x"2b",  x"35", -- 01A0
         x"20",  x"50",  x"4b",  x"54",  x"2e",  x"00",  x"45",  x"49", -- 01A8
         x"4d",  x"45",  x"52",  x"20",  x"49",  x"4d",  x"20",  x"4b", -- 01B0
         x"45",  x"4c",  x"4c",  x"45",  x"52",  x"20",  x"41",  x"55", -- 01B8
         x"53",  x"47",  x"45",  x"53",  x"43",  x"48",  x"2e",  x"3a", -- 01C0
         x"20",  x"2d",  x"78",  x"20",  x"50",  x"4b",  x"54",  x"2e", -- 01C8
         x"20",  x"45",  x"49",  x"4d",  x"45",  x"52",  x"20",  x"5a", -- 01D0
         x"55",  x"4d",  x"20",  x"46",  x"45",  x"4e",  x"53",  x"54", -- 01D8
         x"45",  x"52",  x"20",  x"41",  x"55",  x"53",  x"47",  x"2e", -- 01E0
         x"3a",  x"20",  x"20",  x"20",  x"2b",  x"33",  x"78",  x"20", -- 01E8
         x"50",  x"4b",  x"54",  x"2e",  x"78",  x"20",  x"3d",  x"20", -- 01F0
         x"41",  x"4e",  x"5a",  x"41",  x"48",  x"4c",  x"20",  x"41", -- 01F8
         x"55",  x"46",  x"47",  x"45",  x"46",  x"41",  x"4e",  x"47", -- 0200
         x"2e",  x"20",  x"54",  x"52",  x"4f",  x"50",  x"46",  x"45", -- 0208
         x"4e",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"42", -- 0210
         x"45",  x"49",  x"20",  x"47",  x"55",  x"54",  x"45",  x"4d", -- 0218
         x"20",  x"53",  x"50",  x"49",  x"45",  x"4c",  x"3a",  x"20", -- 0220
         x"20",  x"2b",  x"31",  x"20",  x"53",  x"50",  x"49",  x"45", -- 0228
         x"4c",  x"20",  x"28",  x"4d",  x"41",  x"58",  x"2e",  x"20", -- 0230
         x"33",  x"29",  x"2a",  x"20",  x"45",  x"4e",  x"44",  x"45", -- 0238
         x"20",  x"44",  x"45",  x"53",  x"20",  x"53",  x"50",  x"49", -- 0240
         x"45",  x"4c",  x"45",  x"53",  x"20",  x"2a",  x"cd",  x"00", -- 0248
         x"86",  x"c9",  x"cd",  x"03",  x"86",  x"3a",  x"7f",  x"80", -- 0250
         x"b7",  x"3e",  x"1a",  x"28",  x"0e",  x"dd",  x"2a",  x"7e", -- 0258
         x"80",  x"dd",  x"46",  x"f8",  x"3a",  x"88",  x"80",  x"a0", -- 0260
         x"c0",  x"3e",  x"07",  x"32",  x"0c",  x"80",  x"c9",  x"3e", -- 0268
         x"31",  x"32",  x"7d",  x"80",  x"3e",  x"05",  x"32",  x"63", -- 0270
         x"80",  x"cd",  x"02",  x"92",  x"3a",  x"7d",  x"80",  x"cb", -- 0278
         x"af",  x"32",  x"7d",  x"80",  x"3a",  x"0c",  x"80",  x"b7", -- 0280
         x"28",  x"07",  x"cb",  x"ff",  x"32",  x"0c",  x"80",  x"18", -- 0288
         x"5e",  x"3a",  x"74",  x"80",  x"fe",  x"82",  x"ed",  x"5b", -- 0290
         x"72",  x"80",  x"28",  x"08",  x"11",  x"00",  x"00",  x"3e", -- 0298
         x"13",  x"32",  x"0c",  x"80",  x"3a",  x"80",  x"80",  x"fe", -- 02A0
         x"20",  x"28",  x"05",  x"3e",  x"20",  x"32",  x"0c",  x"80", -- 02A8
         x"ed",  x"53",  x"0d",  x"80",  x"ed",  x"53",  x"86",  x"80", -- 02B0
         x"3e",  x"06",  x"32",  x"88",  x"80",  x"3a",  x"1a",  x"80", -- 02B8
         x"b7",  x"20",  x"2d",  x"3a",  x"c1",  x"81",  x"fe",  x"01", -- 02C0
         x"20",  x"25",  x"e5",  x"d5",  x"11",  x"80",  x"80",  x"21", -- 02C8
         x"07",  x"80",  x"01",  x"05",  x"00",  x"ed",  x"b0",  x"cd", -- 02D0
         x"03",  x"86",  x"dd",  x"2a",  x"7e",  x"80",  x"3e",  x"0a", -- 02D8
         x"d1",  x"ed",  x"53",  x"e1",  x"81",  x"dd",  x"73",  x"fa", -- 02E0
         x"dd",  x"72",  x"f9",  x"dd",  x"77",  x"f8",  x"e1",  x"c9", -- 02E8
         x"01",  x"00",  x"00",  x"ed",  x"43",  x"93",  x"81",  x"3e", -- 02F0
         x"22",  x"32",  x"96",  x"81",  x"ed",  x"53",  x"97",  x"81", -- 02F8
         x"18",  x"ed",  x"7e",  x"fe",  x"0d",  x"28",  x"09",  x"fe", -- 0300
         x"3b",  x"28",  x"05",  x"23",  x"18",  x"f4",  x"18",  x"00", -- 0308
         x"c9",  x"3a",  x"7d",  x"80",  x"cb",  x"ff",  x"18",  x"0c", -- 0310
         x"cd",  x"29",  x"84",  x"7b",  x"32",  x"e4",  x"81",  x"3a", -- 0318
         x"7d",  x"80",  x"cb",  x"f7",  x"32",  x"7d",  x"80",  x"3a", -- 0320
         x"80",  x"80",  x"fe",  x"20",  x"28",  x"05",  x"3e",  x"20", -- 0328
         x"32",  x"0c",  x"80",  x"c9",  x"3a",  x"7d",  x"80",  x"f6", -- 0330
         x"30",  x"32",  x"7d",  x"80",  x"3a",  x"80",  x"80",  x"fe", -- 0338
         x"20",  x"20",  x"07",  x"3e",  x"a1",  x"32",  x"0c",  x"80", -- 0340
         x"18",  x"34",  x"cd",  x"13",  x"a0",  x"3a",  x"0c",  x"80", -- 0348
         x"b7",  x"20",  x"2b",  x"e5",  x"cd",  x"03",  x"86",  x"2a", -- 0350
         x"7e",  x"80",  x"11",  x"00",  x"00",  x"b7",  x"ed",  x"52", -- 0358
         x"3e",  x"06",  x"e5",  x"dd",  x"e1",  x"e1",  x"ca",  x"26", -- 0360
         x"9d",  x"3a",  x"65",  x"a1",  x"b7",  x"ca",  x"4c",  x"9d", -- 0368
         x"ed",  x"5b",  x"72",  x"80",  x"dd",  x"73",  x"fa",  x"dd", -- 0370
         x"72",  x"f9",  x"dd",  x"cb",  x"f8",  x"fe",  x"c3",  x"4c", -- 0378
         x"9d",  x"3a",  x"7d",  x"80",  x"f6",  x"20",  x"32",  x"7d", -- 0380
         x"80",  x"cd",  x"13",  x"a0",  x"3a",  x"6b",  x"a1",  x"3c", -- 0388
         x"32",  x"6b",  x"a1",  x"3a",  x"86",  x"80",  x"32",  x"65", -- 0390
         x"a1",  x"b7",  x"28",  x"11",  x"3a",  x"6b",  x"a1",  x"47", -- 0398
         x"05",  x"3a",  x"6c",  x"a1",  x"3c",  x"b8",  x"20",  x"0d", -- 03A0
         x"32",  x"6c",  x"a1",  x"18",  x"0c",  x"3a",  x"19",  x"80", -- 03A8
         x"cb",  x"87",  x"32",  x"19",  x"80",  x"af",  x"32",  x"65", -- 03B0
         x"a1",  x"3a",  x"80",  x"80",  x"fe",  x"20",  x"28",  x"05", -- 03B8
         x"3e",  x"20",  x"32",  x"0c",  x"80",  x"c3",  x"4c",  x"9d", -- 03C0
         x"3a",  x"6c",  x"a1",  x"47",  x"3a",  x"6b",  x"a1",  x"b7", -- 03C8
         x"28",  x"38",  x"3d",  x"32",  x"6b",  x"a1",  x"4f",  x"3a", -- 03D0
         x"65",  x"a1",  x"b7",  x"79",  x"20",  x"08",  x"3d",  x"b8", -- 03D8
         x"3e",  x"00",  x"20",  x"16",  x"18",  x"0c",  x"b8",  x"3e", -- 03E0
         x"00",  x"20",  x"0f",  x"3a",  x"6c",  x"a1",  x"3d",  x"32", -- 03E8
         x"6c",  x"a1",  x"3a",  x"6d",  x"a1",  x"32",  x"19",  x"80", -- 03F0
         x"3e",  x"01",  x"32",  x"65",  x"a1",  x"3a",  x"80",  x"80"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
