library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom2_4800 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom2_4800;

architecture rtl of rom2_4800 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"82",  x"01",  x"30",  x"d0",  x"88",  x"01",  x"10",  x"00", -- 0000
         x"82",  x"01",  x"30",  x"9c",  x"82",  x"01",  x"10",  x"af", -- 0008
         x"82",  x"01",  x"30",  x"c4",  x"30",  x"c4",  x"84",  x"01", -- 0010
         x"20",  x"9c",  x"82",  x"01",  x"30",  x"83",  x"82",  x"01", -- 0018
         x"20",  x"9c",  x"82",  x"01",  x"08",  x"c4",  x"08",  x"af", -- 0020
         x"82",  x"01",  x"10",  x"9c",  x"82",  x"01",  x"20",  x"af", -- 0028
         x"20",  x"af",  x"00",  x"02",  x"ff",  x"03",  x"80",  x"00", -- 0030
         x"20",  x"e9",  x"82",  x"01",  x"10",  x"dc",  x"82",  x"01", -- 0038
         x"3f",  x"c4",  x"84",  x"01",  x"18",  x"c4",  x"82",  x"01", -- 0040
         x"20",  x"af",  x"82",  x"01",  x"10",  x"9c",  x"82",  x"01", -- 0048
         x"3f",  x"93",  x"00",  x"d5",  x"d6",  x"d7",  x"dd",  x"dc", -- 0050
         x"db",  x"0d",  x"08",  x"07",  x"09",  x"04",  x"08",  x"04", -- 0058
         x"0b",  x"85",  x"fd",  x"88",  x"fd",  x"8b",  x"fd",  x"8e", -- 0060
         x"fd",  x"9a",  x"fd",  x"9d",  x"fd",  x"aa",  x"fd",  x"b6", -- 0068
         x"fd",  x"00",  x"00",  x"00",  x"39",  x"3d",  x"1f",  x"0f", -- 0070
         x"7f",  x"00",  x"00",  x"80",  x"ce",  x"de",  x"fc",  x"f8", -- 0078
         x"ff",  x"ff",  x"0f",  x"1f",  x"3d",  x"39",  x"00",  x"00", -- 0080
         x"00",  x"ff",  x"f8",  x"fc",  x"de",  x"ce",  x"80",  x"00", -- 0088
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"03", -- 0090
         x"07",  x"00",  x"00",  x"00",  x"00",  x"00",  x"80",  x"e0", -- 0098
         x"f0",  x"07",  x"03",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00A0
         x"00",  x"f0",  x"e0",  x"80",  x"00",  x"00",  x"00",  x"00", -- 00A8
         x"00",  x"00",  x"00",  x"00",  x"39",  x"3d",  x"1f",  x"0f", -- 00B0
         x"7f",  x"00",  x"00",  x"80",  x"ce",  x"de",  x"fc",  x"f8", -- 00B8
         x"ff",  x"ff",  x"0f",  x"1f",  x"3d",  x"39",  x"00",  x"00", -- 00C0
         x"00",  x"ff",  x"f8",  x"fc",  x"de",  x"ce",  x"80",  x"00", -- 00C8
         x"00",  x"00",  x"00",  x"00",  x"39",  x"3d",  x"1f",  x"0f", -- 00D0
         x"7f",  x"00",  x"00",  x"80",  x"ce",  x"de",  x"fc",  x"f8", -- 00D8
         x"ff",  x"ff",  x"0f",  x"1f",  x"3d",  x"39",  x"00",  x"00", -- 00E0
         x"00",  x"ff",  x"f8",  x"fc",  x"de",  x"ce",  x"80",  x"00", -- 00E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0100
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0108
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0110
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0118
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0120
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0128
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0130
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0138
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0140
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0148
         x"00",  x"00",  x"70",  x"78",  x"7c",  x"3e",  x"3e",  x"3e", -- 0150
         x"1e",  x"00",  x"07",  x"0f",  x"1f",  x"3e",  x"3e",  x"3e", -- 0158
         x"3c",  x"1e",  x"1e",  x"3e",  x"3e",  x"3c",  x"18",  x"00", -- 0160
         x"00",  x"3c",  x"3c",  x"3e",  x"3f",  x"1f",  x"0c",  x"00", -- 0168
         x"00",  x"00",  x"70",  x"78",  x"7c",  x"3e",  x"3e",  x"3e", -- 0170
         x"1e",  x"00",  x"07",  x"0f",  x"1f",  x"3e",  x"3e",  x"3e", -- 0178
         x"3c",  x"1e",  x"1e",  x"3e",  x"3e",  x"3c",  x"18",  x"00", -- 0180
         x"00",  x"3c",  x"3c",  x"3e",  x"3f",  x"1f",  x"0c",  x"00", -- 0188
         x"00",  x"00",  x"70",  x"78",  x"7c",  x"3e",  x"3e",  x"3e", -- 0190
         x"1e",  x"00",  x"07",  x"0f",  x"1f",  x"3e",  x"3e",  x"3e", -- 0198
         x"3c",  x"1e",  x"1e",  x"3e",  x"3e",  x"3c",  x"18",  x"00", -- 01A0
         x"00",  x"3c",  x"3c",  x"3e",  x"3f",  x"1f",  x"0c",  x"00", -- 01A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01C8
         x"00",  x"00",  x"00",  x"30",  x"38",  x"1c",  x"00",  x"00", -- 01D0
         x"00",  x"00",  x"00",  x"06",  x"0e",  x"1c",  x"00",  x"00", -- 01D8
         x"00",  x"04",  x"0e",  x"16",  x"38",  x"18",  x"00",  x"00", -- 01E0
         x"00",  x"10",  x"38",  x"34",  x"0e",  x"0c",  x"00",  x"00", -- 01E8
         x"00",  x"00",  x"50",  x"30",  x"7c",  x"1c",  x"21",  x"30", -- 01F0
         x"11",  x"00",  x"05",  x"06",  x"1f",  x"1c",  x"42",  x"06", -- 01F8
         x"44",  x"04",  x"1f",  x"16",  x"7d",  x"38",  x"08",  x"00", -- 0200
         x"00",  x"10",  x"7c",  x"34",  x"5f",  x"0e",  x"08",  x"00", -- 0208
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0210
         x"00",  x"00",  x"00",  x"00",  x"06",  x"14",  x"18",  x"00", -- 0218
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0220
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0228
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0230
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0238
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0240
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0248
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0250
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0258
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0260
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0268
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0270
         x"00",  x"00",  x"00",  x"00",  x"60",  x"28",  x"18",  x"00", -- 0278
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0280
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0288
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0290
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0298
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02C8
         x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02D0
         x"00",  x"3f",  x"3f",  x"3f",  x"3f",  x"3f",  x"3f",  x"3f", -- 02D8
         x"00",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f", -- 02E0
         x"00",  x"03",  x"03",  x"03",  x"03",  x"03",  x"03",  x"03", -- 02E8
         x"7f",  x"02",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02F0
         x"00",  x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 02F8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"c6",  x"c2",  x"e0", -- 0300
         x"f3",  x"87",  x"ff",  x"ff",  x"7f",  x"31",  x"21",  x"83", -- 0308
         x"e7",  x"f0",  x"07",  x"f3",  x"e0",  x"c2",  x"c6",  x"ff", -- 0310
         x"ff",  x"ff",  x"f0",  x"e7",  x"83",  x"21",  x"31",  x"7f", -- 0318
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"c6",  x"c2",  x"e0", -- 0320
         x"f3",  x"87",  x"ff",  x"ff",  x"7f",  x"31",  x"21",  x"83", -- 0328
         x"e7",  x"f0",  x"07",  x"f3",  x"e0",  x"c2",  x"c6",  x"ff", -- 0330
         x"ff",  x"ff",  x"f0",  x"e7",  x"83",  x"21",  x"31",  x"7f", -- 0338
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"c6",  x"c2",  x"e0", -- 0340
         x"f3",  x"87",  x"ff",  x"ff",  x"7f",  x"31",  x"21",  x"83", -- 0348
         x"e7",  x"f0",  x"07",  x"f3",  x"e0",  x"c2",  x"c6",  x"ff", -- 0350
         x"ff",  x"ff",  x"f0",  x"e7",  x"83",  x"21",  x"31",  x"7f", -- 0358
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0360
         x"fc",  x"f8",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f", -- 0368
         x"1f",  x"0f",  x"f8",  x"fc",  x"ff",  x"ff",  x"ff",  x"ff", -- 0370
         x"ff",  x"ff",  x"0f",  x"1f",  x"7f",  x"ff",  x"ff",  x"ff", -- 0378
         x"ff",  x"ff",  x"f3",  x"fd",  x"fe",  x"fe",  x"fe",  x"fe", -- 0380
         x"fe",  x"fe",  x"e7",  x"5f",  x"3f",  x"3f",  x"3f",  x"3f", -- 0388
         x"3f",  x"3f",  x"fe",  x"fe",  x"fe",  x"fe",  x"ff",  x"ff", -- 0390
         x"ff",  x"ff",  x"3f",  x"3f",  x"3f",  x"3f",  x"7f",  x"7f", -- 0398
         x"ff",  x"ff",  x"f3",  x"8d",  x"86",  x"82",  x"c0",  x"c0", -- 03A0
         x"c0",  x"e0",  x"e7",  x"58",  x"30",  x"20",  x"01",  x"01", -- 03A8
         x"01",  x"03",  x"e0",  x"e0",  x"c0",  x"80",  x"83",  x"e7", -- 03B0
         x"ff",  x"ff",  x"03",  x"03",  x"01",  x"00",  x"60",  x"73", -- 03B8
         x"ff",  x"ff",  x"f3",  x"8d",  x"86",  x"82",  x"c0",  x"c0", -- 03C0
         x"c0",  x"e0",  x"e7",  x"58",  x"30",  x"20",  x"01",  x"01", -- 03C8
         x"01",  x"03",  x"e0",  x"e0",  x"c0",  x"80",  x"83",  x"e7", -- 03D0
         x"ff",  x"ff",  x"03",  x"03",  x"01",  x"00",  x"60",  x"73", -- 03D8
         x"ff",  x"ff",  x"f3",  x"8d",  x"86",  x"82",  x"c0",  x"c0", -- 03E0
         x"c0",  x"e0",  x"e7",  x"58",  x"30",  x"20",  x"01",  x"01", -- 03E8
         x"01",  x"03",  x"e0",  x"e0",  x"c0",  x"80",  x"83",  x"e7", -- 03F0
         x"ff",  x"ff",  x"03",  x"03",  x"01",  x"00",  x"60",  x"73"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
