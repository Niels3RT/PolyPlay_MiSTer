library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_zre_0400 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_zre_0400;

architecture rtl of rom_zre_0400 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"b7",  x"21",  x"16",  x"00",  x"fd",  x"cb",  x"00",  x"46", -- 0000
         x"20",  x"03",  x"21",  x"0e",  x"00",  x"ed",  x"42",  x"da", -- 0008
         x"97",  x"05",  x"20",  x"14",  x"21",  x"09",  x"0d",  x"36", -- 0010
         x"01",  x"cd",  x"73",  x"06",  x"3a",  x"1a",  x"0d",  x"47", -- 0018
         x"2a",  x"01",  x"0d",  x"23",  x"36",  x"80",  x"10",  x"fb", -- 0020
         x"cd",  x"37",  x"04",  x"2a",  x"01",  x"0d",  x"cd",  x"73", -- 0028
         x"06",  x"21",  x"09",  x"0d",  x"36",  x"2f",  x"c9",  x"11", -- 0030
         x"c0",  x"f8",  x"21",  x"00",  x"f9",  x"01",  x"c0",  x"00", -- 0038
         x"ed",  x"b0",  x"cd",  x"22",  x"06",  x"01",  x"40",  x"01", -- 0040
         x"ed",  x"b0",  x"e5",  x"d5",  x"fd",  x"cb",  x"00",  x"46", -- 0048
         x"20",  x"20",  x"21",  x"05",  x"0d",  x"3a",  x"03",  x"0d", -- 0050
         x"77",  x"3a",  x"55",  x"0d",  x"47",  x"3a",  x"00",  x"0d", -- 0058
         x"cb",  x"2f",  x"c6",  x"de",  x"b8",  x"30",  x"03",  x"34", -- 0060
         x"18",  x"15",  x"d6",  x"08",  x"b8",  x"38",  x"10",  x"35", -- 0068
         x"18",  x"0d",  x"db",  x"84",  x"1f",  x"1f",  x"f5",  x"d4", -- 0070
         x"cd",  x"05",  x"f1",  x"1f",  x"d4",  x"e4",  x"05",  x"21", -- 0078
         x"a0",  x"fa",  x"3a",  x"00",  x"0d",  x"47",  x"3a",  x"05", -- 0080
         x"0d",  x"80",  x"fe",  x"40",  x"38",  x"04",  x"fe",  x"c0", -- 0088
         x"38",  x"5d",  x"32",  x"00",  x"0d",  x"cb",  x"2f",  x"85", -- 0090
         x"6f",  x"3e",  x"80",  x"be",  x"38",  x"4c",  x"11",  x"a5", -- 0098
         x"13",  x"3a",  x"05",  x"0d",  x"c6",  x"04",  x"83",  x"5f", -- 00A0
         x"30",  x"01",  x"14",  x"1a",  x"06",  x"03",  x"2b",  x"4f", -- 00A8
         x"3e",  x"7f",  x"be",  x"38",  x"01",  x"71",  x"23",  x"0c", -- 00B0
         x"10",  x"f8",  x"d1",  x"e1",  x"cd",  x"d8",  x"06",  x"cd", -- 00B8
         x"22",  x"06",  x"01",  x"00",  x"05",  x"fd",  x"cb",  x"00", -- 00C0
         x"46",  x"20",  x"03",  x"01",  x"00",  x"03",  x"ed",  x"b0", -- 00C8
         x"c9",  x"c5",  x"11",  x"c0",  x"f8",  x"21",  x"00",  x"f9", -- 00D0
         x"01",  x"00",  x"07",  x"fd",  x"cb",  x"00",  x"46",  x"20", -- 00D8
         x"03",  x"01",  x"00",  x"05",  x"ed",  x"b0",  x"c1",  x"10", -- 00E0
         x"e8",  x"c9",  x"3e",  x"9e",  x"be",  x"20",  x"5e",  x"fd", -- 00E8
         x"cb",  x"00",  x"46",  x"28",  x"58",  x"21",  x"49",  x"15", -- 00F0
         x"cd",  x"e0",  x"01",  x"d1",  x"e1",  x"01",  x"40",  x"00", -- 00F8
         x"ed",  x"b0",  x"21",  x"c0",  x"fa",  x"22",  x"1b",  x"0d", -- 0100
         x"3a",  x"05",  x"0d",  x"cb",  x"7f",  x"16",  x"01",  x"28", -- 0108
         x"08",  x"16",  x"ff",  x"21",  x"fa",  x"fa",  x"22",  x"1b", -- 0110
         x"0d",  x"06",  x"05",  x"0e",  x"80",  x"18",  x"02",  x"0e", -- 0118
         x"af",  x"cd",  x"33",  x"07",  x"0d",  x"3e",  x"50",  x"b9", -- 0120
         x"20",  x"f7",  x"21",  x"00",  x"08",  x"2b",  x"7d",  x"b4", -- 0128
         x"20",  x"fb",  x"0e",  x"50",  x"cd",  x"33",  x"07",  x"0c", -- 0130
         x"3e",  x"01",  x"b8",  x"3e",  x"af",  x"20",  x"02",  x"3e", -- 0138
         x"ff",  x"b9",  x"20",  x"f0",  x"10",  x"d9",  x"0e",  x"01", -- 0140
         x"cd",  x"33",  x"07",  x"18",  x"16",  x"cd",  x"22",  x"06", -- 0148
         x"d1",  x"e1",  x"01",  x"40",  x"00",  x"ed",  x"b0",  x"fd", -- 0150
         x"cb",  x"00",  x"46",  x"28",  x"06",  x"21",  x"50",  x"15", -- 0158
         x"cd",  x"d4",  x"01",  x"f1",  x"cd",  x"f0",  x"05",  x"61", -- 0160
         x"14",  x"21",  x"6a",  x"f9",  x"22",  x"3f",  x"0c",  x"21", -- 0168
         x"2c",  x"01",  x"f1",  x"c1",  x"b7",  x"ed",  x"42",  x"22", -- 0170
         x"3d",  x"0c",  x"cd",  x"70",  x"02",  x"cd",  x"f0",  x"05", -- 0178
         x"7d",  x"14",  x"21",  x"1a",  x"0d",  x"7e",  x"dd",  x"77", -- 0180
         x"00",  x"cb",  x"2f",  x"86",  x"fe",  x"20",  x"36",  x"1e", -- 0188
         x"d2",  x"85",  x"12",  x"77",  x"c3",  x"85",  x"12",  x"cd", -- 0190
         x"37",  x"04",  x"21",  x"04",  x"0d",  x"35",  x"20",  x"08", -- 0198
         x"36",  x"07",  x"cd",  x"c5",  x"05",  x"32",  x"03",  x"0d", -- 01A0
         x"2a",  x"01",  x"0d",  x"3a",  x"03",  x"0d",  x"85",  x"fe", -- 01A8
         x"c0",  x"28",  x"0e",  x"47",  x"3a",  x"1a",  x"0d",  x"80", -- 01B0
         x"fe",  x"fe",  x"78",  x"28",  x"04",  x"6f",  x"22",  x"01", -- 01B8
         x"0d",  x"cd",  x"73",  x"06",  x"c9",  x"ed",  x"5f",  x"e6", -- 01C0
         x"03",  x"c8",  x"3d",  x"3d",  x"c9",  x"3a",  x"05",  x"0d", -- 01C8
         x"3c",  x"fa",  x"d7",  x"05",  x"fe",  x"05",  x"d0",  x"32", -- 01D0
         x"05",  x"0d",  x"21",  x"56",  x"0c",  x"3e",  x"90",  x"be", -- 01D8
         x"d8",  x"34",  x"34",  x"c9",  x"3a",  x"05",  x"0d",  x"3d", -- 01E0
         x"f2",  x"d7",  x"05",  x"fe",  x"fc",  x"d8",  x"18",  x"e7", -- 01E8
         x"e1",  x"5e",  x"23",  x"56",  x"23",  x"e5",  x"d5",  x"e1", -- 01F0
         x"5e",  x"23",  x"56",  x"23",  x"4e",  x"06",  x"00",  x"23", -- 01F8
         x"ed",  x"b0",  x"c9",  x"3e",  x"4d",  x"32",  x"bf",  x"0c", -- 0200
         x"fd",  x"cb",  x"00",  x"46",  x"20",  x"0b",  x"c5",  x"cd", -- 0208
         x"9a",  x"01",  x"c1",  x"c0",  x"3a",  x"03",  x"0c",  x"b7", -- 0210
         x"c0",  x"3a",  x"bf",  x"0c",  x"b7",  x"20",  x"e9",  x"10", -- 0218
         x"e2",  x"c9",  x"d5",  x"e5",  x"21",  x"a0",  x"fa",  x"3a", -- 0220
         x"00",  x"0d",  x"cb",  x"2f",  x"85",  x"6f",  x"c5",  x"01", -- 0228
         x"3f",  x"ff",  x"09",  x"11",  x"0a",  x"0d",  x"06",  x"03", -- 0230
         x"cd",  x"69",  x"06",  x"01",  x"3c",  x"00",  x"09",  x"06", -- 0238
         x"05",  x"cd",  x"69",  x"06",  x"01",  x"3b",  x"00",  x"09", -- 0240
         x"06",  x"05",  x"cd",  x"69",  x"06",  x"01",  x"3c",  x"00", -- 0248
         x"09",  x"06",  x"03",  x"cd",  x"69",  x"06",  x"c1",  x"e1", -- 0250
         x"d1",  x"c9",  x"d5",  x"e5",  x"21",  x"a0",  x"ff",  x"fd", -- 0258
         x"cb",  x"00",  x"46",  x"20",  x"c9",  x"25",  x"25",  x"18", -- 0260
         x"c5",  x"1a",  x"4e",  x"77",  x"79",  x"12",  x"23",  x"13", -- 0268
         x"10",  x"f7",  x"c9",  x"21",  x"09",  x"0d",  x"35",  x"fa", -- 0270
         x"be",  x"06",  x"28",  x"01",  x"c9",  x"21",  x"c0",  x"ff", -- 0278
         x"fd",  x"cb",  x"00",  x"46",  x"20",  x"08",  x"3a",  x"01", -- 0280
         x"0d",  x"32",  x"55",  x"0d",  x"25",  x"25",  x"3a",  x"01", -- 0288
         x"0d",  x"95",  x"3d",  x"28",  x"06",  x"47",  x"23",  x"36", -- 0290
         x"91",  x"10",  x"fb",  x"23",  x"3a",  x"08",  x"0d",  x"ee", -- 0298
         x"03",  x"32",  x"08",  x"0d",  x"77",  x"e5",  x"21",  x"1a", -- 02A0
         x"0d",  x"46",  x"e1",  x"23",  x"36",  x"20",  x"10",  x"fb", -- 02A8
         x"23",  x"77",  x"3e",  x"ff",  x"95",  x"3d",  x"c8",  x"47", -- 02B0
         x"23",  x"36",  x"91",  x"10",  x"fb",  x"c9",  x"36",  x"0f", -- 02B8
         x"21",  x"c0",  x"ff",  x"fd",  x"cb",  x"00",  x"46",  x"20", -- 02C0
         x"02",  x"25",  x"25",  x"36",  x"9e",  x"06",  x"3f",  x"3e", -- 02C8
         x"20",  x"23",  x"77",  x"10",  x"fc",  x"36",  x"9e",  x"c9", -- 02D0
         x"e5",  x"c5",  x"0e",  x"ba",  x"3a",  x"05",  x"0d",  x"cb", -- 02D8
         x"7f",  x"20",  x"01",  x"3c",  x"cb",  x"2f",  x"47",  x"cb", -- 02E0
         x"27",  x"cb",  x"27",  x"80",  x"cb",  x"27",  x"81",  x"4f", -- 02E8
         x"21",  x"0a",  x"0d",  x"3e",  x"a0",  x"06",  x"03",  x"77", -- 02F0
         x"3c",  x"23",  x"10",  x"fb",  x"71",  x"23",  x"0c",  x"06", -- 02F8
         x"03",  x"77",  x"3c",  x"23",  x"10",  x"fb",  x"06",  x"09", -- 0300
         x"71",  x"23",  x"0c",  x"10",  x"fb",  x"c1",  x"e1",  x"c9", -- 0308
         x"e5",  x"c5",  x"36",  x"20",  x"3e",  x"d8",  x"06",  x"04", -- 0310
         x"23",  x"77",  x"3c",  x"10",  x"fb",  x"23",  x"36",  x"20", -- 0318
         x"01",  x"3b",  x"00",  x"09",  x"36",  x"20",  x"06",  x"04", -- 0320
         x"23",  x"77",  x"3c",  x"10",  x"fb",  x"23",  x"36",  x"20", -- 0328
         x"c1",  x"e1",  x"c9",  x"3e",  x"05",  x"d3",  x"80",  x"79", -- 0330
         x"d3",  x"80",  x"1e",  x"06",  x"79",  x"e6",  x"0f",  x"20", -- 0338
         x"0c",  x"2a",  x"1b",  x"0d",  x"7d",  x"82",  x"6f",  x"22", -- 0340
         x"1b",  x"0d",  x"cd",  x"10",  x"07",  x"79",  x"2f",  x"3d", -- 0348
         x"20",  x"fd",  x"1d",  x"20",  x"f8",  x"c9",  x"e5",  x"c5", -- 0350
         x"06",  x"3a",  x"3e",  x"9f",  x"cd",  x"8b",  x"07",  x"c1", -- 0358
         x"e1",  x"c9",  x"e5",  x"c5",  x"36",  x"9f",  x"23",  x"3e", -- 0360
         x"20",  x"06",  x"06",  x"cd",  x"8b",  x"07",  x"36",  x"9f", -- 0368
         x"23",  x"06",  x"0e",  x"cd",  x"8b",  x"07",  x"36",  x"9f", -- 0370
         x"23",  x"06",  x"12",  x"cd",  x"8b",  x"07",  x"36",  x"9f", -- 0378
         x"23",  x"06",  x"0f",  x"cd",  x"8b",  x"07",  x"36",  x"9f", -- 0380
         x"c1",  x"e1",  x"c9",  x"77",  x"23",  x"10",  x"fc",  x"c9", -- 0388
         x"eb",  x"c5",  x"4e",  x"23",  x"06",  x"00",  x"ed",  x"b0", -- 0390
         x"eb",  x"c1",  x"c9",  x"cb",  x"27",  x"32",  x"3d",  x"0c", -- 0398
         x"cd",  x"70",  x"02",  x"2b",  x"2b",  x"2b",  x"7e",  x"36", -- 03A0
         x"2c",  x"23",  x"77",  x"23",  x"11",  x"1d",  x"15",  x"cd", -- 03A8
         x"90",  x"07",  x"c9",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
