library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom2_2000 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom2_2000;

architecture rtl of rom2_2000 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"46",  x"0c",  x"ed",  x"b0",  x"3e",  x"05",  x"32",  x"c1", -- 0000
         x"0c",  x"cd",  x"2e",  x"20",  x"c9",  x"21",  x"4a",  x"0c", -- 0008
         x"73",  x"f5",  x"2a",  x"48",  x"0c",  x"7d",  x"81",  x"e6", -- 0010
         x"3f",  x"fe",  x"3f",  x"30",  x"0f",  x"6f",  x"7c",  x"80", -- 0018
         x"e6",  x"1f",  x"28",  x"08",  x"fe",  x"1f",  x"30",  x"04", -- 0020
         x"67",  x"22",  x"48",  x"0c",  x"f1",  x"c9",  x"11",  x"a3", -- 0028
         x"23",  x"3a",  x"b2",  x"0c",  x"e6",  x"03",  x"87",  x"87", -- 0030
         x"83",  x"5f",  x"30",  x"01",  x"14",  x"2a",  x"ae",  x"0c", -- 0038
         x"01",  x"3f",  x"00",  x"cd",  x"88",  x"1f",  x"09",  x"cd", -- 0040
         x"88",  x"1f",  x"c9",  x"af",  x"2a",  x"ae",  x"0c",  x"01", -- 0048
         x"3f",  x"00",  x"cd",  x"5c",  x"1f",  x"09",  x"cd",  x"5c", -- 0050
         x"1f",  x"c9",  x"2a",  x"46",  x"0c",  x"01",  x"3f",  x"00", -- 0058
         x"af",  x"cd",  x"a8",  x"1f",  x"c0",  x"09",  x"cd",  x"a8", -- 0060
         x"1f",  x"c9",  x"2a",  x"48",  x"0c",  x"cb",  x"05",  x"cb", -- 0068
         x"05",  x"cb",  x"3c",  x"cb",  x"1d",  x"cb",  x"3c",  x"cb", -- 0070
         x"1d",  x"11",  x"00",  x"f8",  x"19",  x"22",  x"46",  x"0c", -- 0078
         x"c9",  x"21",  x"b8",  x"0c",  x"7e",  x"b7",  x"c8",  x"35", -- 0080
         x"20",  x"06",  x"2a",  x"b3",  x"0c",  x"36",  x"00",  x"c9", -- 0088
         x"3a",  x"b7",  x"0c",  x"e6",  x"03",  x"87",  x"21",  x"b0", -- 0090
         x"23",  x"85",  x"6f",  x"30",  x"01",  x"24",  x"5e",  x"23", -- 0098
         x"56",  x"2a",  x"b5",  x"0c",  x"7d",  x"83",  x"cb",  x"77", -- 00A0
         x"20",  x"41",  x"e6",  x"3f",  x"6f",  x"7c",  x"82",  x"e6", -- 00A8
         x"1f",  x"fe",  x"01",  x"38",  x"36",  x"67",  x"22",  x"48", -- 00B0
         x"0c",  x"cd",  x"6a",  x"20",  x"2a",  x"b3",  x"0c",  x"7e", -- 00B8
         x"fe",  x"b5",  x"20",  x"02",  x"36",  x"00",  x"2a",  x"46", -- 00C0
         x"0c",  x"7e",  x"b7",  x"28",  x"0b",  x"21",  x"b8",  x"0c", -- 00C8
         x"36",  x"00",  x"fe",  x"ab",  x"c8",  x"fe",  x"ac",  x"c8", -- 00D0
         x"21",  x"46",  x"0c",  x"11",  x"b3",  x"0c",  x"01",  x"04", -- 00D8
         x"00",  x"ed",  x"b0",  x"2a",  x"b3",  x"0c",  x"3e",  x"b5", -- 00E0
         x"77",  x"b7",  x"c9",  x"2a",  x"b3",  x"0c",  x"7e",  x"fe", -- 00E8
         x"b5",  x"20",  x"02",  x"36",  x"00",  x"af",  x"32",  x"b8", -- 00F0
         x"0c",  x"c9",  x"21",  x"c3",  x"0c",  x"7e",  x"b7",  x"c0", -- 00F8
         x"db",  x"84",  x"ee",  x"00",  x"cb",  x"47",  x"c0",  x"3e", -- 0100
         x"14",  x"32",  x"c3",  x"0c",  x"21",  x"b0",  x"0c",  x"11", -- 0108
         x"b5",  x"0c",  x"01",  x"03",  x"00",  x"ed",  x"b0",  x"3a", -- 0110
         x"b7",  x"0c",  x"cb",  x"4f",  x"3e",  x"14",  x"28",  x"02", -- 0118
         x"cb",  x"3f",  x"12",  x"21",  x"b5",  x"0c",  x"3a",  x"b7", -- 0120
         x"0c",  x"fe",  x"01",  x"28",  x"07",  x"34",  x"23",  x"fe", -- 0128
         x"03",  x"38",  x"01",  x"34",  x"cd",  x"90",  x"20",  x"c8", -- 0130
         x"21",  x"1c",  x"0c",  x"35",  x"af",  x"32",  x"bf",  x"0c", -- 0138
         x"3e",  x"0a",  x"3c",  x"32",  x"c0",  x"0c",  x"c9",  x"21", -- 0140
         x"00",  x"f8",  x"11",  x"0a",  x"00",  x"19",  x"22",  x"3f", -- 0148
         x"0c",  x"2a",  x"06",  x"0c",  x"22",  x"3d",  x"0c",  x"cd", -- 0150
         x"70",  x"02",  x"21",  x"00",  x"f8",  x"11",  x"1b",  x"00", -- 0158
         x"19",  x"22",  x"3f",  x"0c",  x"2a",  x"18",  x"0c",  x"22", -- 0160
         x"3d",  x"0c",  x"cd",  x"70",  x"02",  x"21",  x"00",  x"f8", -- 0168
         x"11",  x"3b",  x"00",  x"19",  x"22",  x"3f",  x"0c",  x"2a", -- 0170
         x"1c",  x"0c",  x"22",  x"3d",  x"0c",  x"cd",  x"70",  x"02", -- 0178
         x"3a",  x"bf",  x"0c",  x"b7",  x"c0",  x"3a",  x"c0",  x"0c", -- 0180
         x"3d",  x"20",  x"27",  x"21",  x"c0",  x"23",  x"cd",  x"d4", -- 0188
         x"01",  x"3a",  x"c4",  x"0c",  x"3d",  x"32",  x"c4",  x"0c", -- 0190
         x"20",  x"09",  x"21",  x"c0",  x"0c",  x"35",  x"3e",  x"19", -- 0198
         x"32",  x"c4",  x"0c",  x"3e",  x"0a",  x"32",  x"bf",  x"0c", -- 01A0
         x"21",  x"00",  x"f8",  x"11",  x"2d",  x"00",  x"19",  x"36", -- 01A8
         x"92",  x"c9",  x"fe",  x"f0",  x"30",  x"0b",  x"32",  x"c0", -- 01B0
         x"0c",  x"21",  x"c0",  x"23",  x"cd",  x"d4",  x"01",  x"18", -- 01B8
         x"13",  x"21",  x"1c",  x"0c",  x"7e",  x"b7",  x"28",  x"0c", -- 01C0
         x"35",  x"3e",  x"0a",  x"32",  x"c0",  x"0c",  x"21",  x"66", -- 01C8
         x"24",  x"cd",  x"d4",  x"01",  x"3e",  x"4b",  x"32",  x"bf", -- 01D0
         x"0c",  x"21",  x"00",  x"f8",  x"11",  x"2d",  x"00",  x"19", -- 01D8
         x"3a",  x"c0",  x"0c",  x"3d",  x"cb",  x"7f",  x"20",  x"05", -- 01E0
         x"36",  x"91",  x"2b",  x"18",  x"f6",  x"36",  x"00",  x"c9", -- 01E8
         x"3d",  x"3d",  x"20",  x"52",  x"45",  x"43",  x"4f",  x"52", -- 01F0
         x"44",  x"3a",  x"30",  x"30",  x"20",  x"3d",  x"3d",  x"3d", -- 01F8
         x"3d",  x"3d",  x"20",  x"54",  x"52",  x"45",  x"46",  x"46", -- 0200
         x"45",  x"52",  x"3a",  x"30",  x"30",  x"20",  x"3d",  x"3d", -- 0208
         x"3d",  x"3d",  x"3d",  x"20",  x"00",  x"00",  x"00",  x"00", -- 0210
         x"00",  x"00",  x"00",  x"00",  x"00",  x"0f",  x"00",  x"3d", -- 0218
         x"3d",  x"3d",  x"3d",  x"20",  x"53",  x"43",  x"48",  x"55", -- 0220
         x"53",  x"53",  x"3a",  x"30",  x"30",  x"20",  x"3d",  x"3d", -- 0228
         x"20",  x"4b",  x"45",  x"49",  x"4e",  x"45",  x"4e",  x"20", -- 0230
         x"53",  x"43",  x"48",  x"55",  x"53",  x"53",  x"20",  x"4d", -- 0238
         x"45",  x"48",  x"52",  x"20",  x"2d",  x"20",  x"45",  x"4e", -- 0240
         x"44",  x"45",  x"20",  x"44",  x"45",  x"53",  x"20",  x"53", -- 0248
         x"50",  x"49",  x"45",  x"4c",  x"45",  x"53",  x"20",  x"44", -- 0250
         x"45",  x"52",  x"20",  x"44",  x"41",  x"56",  x"4f",  x"4e", -- 0258
         x"4c",  x"41",  x"55",  x"46",  x"45",  x"4e",  x"44",  x"45", -- 0260
         x"20",  x"48",  x"49",  x"52",  x"53",  x"43",  x"48",  x"20", -- 0268
         x"53",  x"4f",  x"4c",  x"4c",  x"20",  x"56",  x"45",  x"52", -- 0270
         x"46",  x"4f",  x"4c",  x"47",  x"54",  x"20",  x"55",  x"4e", -- 0278
         x"44",  x"20",  x"45",  x"52",  x"4c",  x"45",  x"47",  x"54", -- 0280
         x"20",  x"57",  x"45",  x"52",  x"44",  x"45",  x"4e",  x"2e", -- 0288
         x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"44", -- 0290
         x"41",  x"46",  x"55",  x"45",  x"52",  x"20",  x"53",  x"54", -- 0298
         x"45",  x"48",  x"45",  x"4e",  x"20",  x"31",  x"30",  x"20", -- 02A0
         x"53",  x"43",  x"48",  x"55",  x"53",  x"53",  x"20",  x"5a", -- 02A8
         x"55",  x"52",  x"20",  x"56",  x"45",  x"52",  x"46",  x"55", -- 02B0
         x"45",  x"47",  x"55",  x"4e",  x"47",  x"2e",  x"45",  x"49", -- 02B8
         x"4e",  x"20",  x"53",  x"43",  x"48",  x"55",  x"53",  x"53", -- 02C0
         x"2c",  x"44",  x"45",  x"52",  x"20",  x"44",  x"45",  x"4e", -- 02C8
         x"20",  x"48",  x"49",  x"52",  x"53",  x"43",  x"48",  x"20", -- 02D0
         x"54",  x"52",  x"49",  x"46",  x"46",  x"54",  x"2c",  x"57", -- 02D8
         x"49",  x"52",  x"44",  x"20",  x"4e",  x"49",  x"43",  x"48", -- 02E0
         x"54",  x"20",  x"41",  x"42",  x"47",  x"45",  x"5a",  x"4f", -- 02E8
         x"47",  x"45",  x"4e",  x"2e",  x"45",  x"54",  x"57",  x"41", -- 02F0
         x"20",  x"41",  x"4c",  x"4c",  x"45",  x"52",  x"20",  x"31", -- 02F8
         x"35",  x"20",  x"53",  x"45",  x"4b",  x"55",  x"4e",  x"44", -- 0300
         x"45",  x"4e",  x"20",  x"4d",  x"55",  x"53",  x"53",  x"20", -- 0308
         x"45",  x"49",  x"4e",  x"20",  x"53",  x"43",  x"48",  x"55", -- 0310
         x"53",  x"53",  x"20",  x"41",  x"42",  x"47",  x"45",  x"47", -- 0318
         x"45",  x"42",  x"45",  x"4e",  x"20",  x"57",  x"45",  x"52", -- 0320
         x"44",  x"45",  x"4e",  x"2c",  x"53",  x"4f",  x"4e",  x"53", -- 0328
         x"54",  x"20",  x"47",  x"45",  x"48",  x"54",  x"20",  x"44", -- 0330
         x"49",  x"45",  x"53",  x"45",  x"52",  x"20",  x"53",  x"43", -- 0338
         x"48",  x"55",  x"53",  x"53",  x"20",  x"56",  x"45",  x"52", -- 0340
         x"4c",  x"4f",  x"52",  x"45",  x"4e",  x"2e",  x"57",  x"45", -- 0348
         x"49",  x"44",  x"4d",  x"41",  x"4e",  x"4e",  x"53",  x"20", -- 0350
         x"48",  x"45",  x"49",  x"4c",  x"20",  x"21",  x"30",  x"01", -- 0358
         x"88",  x"01",  x"1e",  x"02",  x"35",  x"03",  x"0f",  x"04", -- 0360
         x"2c",  x"05",  x"06",  x"06",  x"bb",  x"06",  x"e2",  x"06", -- 0368
         x"e0",  x"f8",  x"20",  x"03",  x"03",  x"05",  x"93",  x"94", -- 0370
         x"95",  x"96",  x"97",  x"98",  x"99",  x"9a",  x"9b",  x"9f", -- 0378
         x"a0",  x"a1",  x"a2",  x"a3",  x"a4",  x"a5",  x"a6",  x"a7", -- 0380
         x"93",  x"94",  x"95",  x"96",  x"97",  x"98",  x"9c",  x"9d", -- 0388
         x"9e",  x"9f",  x"a0",  x"a1",  x"a2",  x"a3",  x"a4",  x"a8", -- 0390
         x"a9",  x"aa",  x"00",  x"00",  x"00",  x"b6",  x"b7",  x"b8", -- 0398
         x"b9",  x"ba",  x"bb",  x"ad",  x"ae",  x"af",  x"b0",  x"b1", -- 03A0
         x"b2",  x"b3",  x"b4",  x"20",  x"04",  x"20",  x"10",  x"00", -- 03A8
         x"01",  x"00",  x"ff",  x"00",  x"00",  x"ff",  x"00",  x"01", -- 03B0
         x"01",  x"ff",  x"ff",  x"ff",  x"01",  x"01",  x"ff",  x"01", -- 03B8
         x"03",  x"30",  x"00",  x"50",  x"12",  x"82",  x"01",  x"18", -- 03C0
         x"dc",  x"82",  x"01",  x"08",  x"af",  x"82",  x"01",  x"10", -- 03C8
         x"af",  x"82",  x"01",  x"10",  x"af",  x"82",  x"01",  x"30", -- 03D0
         x"af",  x"82",  x"01",  x"10",  x"93",  x"82",  x"01",  x"10", -- 03D8
         x"93",  x"82",  x"01",  x"10",  x"a5",  x"82",  x"01",  x"10", -- 03E0
         x"a5",  x"82",  x"01",  x"10",  x"af",  x"82",  x"01",  x"18", -- 03E8
         x"af",  x"82",  x"01",  x"08",  x"c4",  x"82",  x"01",  x"10", -- 03F0
         x"c4",  x"82",  x"01",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
