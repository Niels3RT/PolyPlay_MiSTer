library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom2_2800 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom2_2800;

architecture rtl of rom2_2800 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"21",  x"18",  x"0c",  x"11",  x"19",  x"0c",  x"01",  x"c8", -- 0000
         x"00",  x"36",  x"00",  x"ed",  x"b0",  x"cd",  x"b7",  x"02", -- 0008
         x"21",  x"62",  x"00",  x"11",  x"db",  x"3c",  x"01",  x"f0", -- 0010
         x"00",  x"cd",  x"c8",  x"02",  x"21",  x"5e",  x"00",  x"11", -- 0018
         x"cb",  x"3d",  x"01",  x"90",  x"00",  x"cd",  x"ce",  x"02", -- 0020
         x"21",  x"5e",  x"00",  x"11",  x"5b",  x"3e",  x"01",  x"d0", -- 0028
         x"00",  x"cd",  x"d4",  x"02",  x"cd",  x"97",  x"2e",  x"21", -- 0030
         x"84",  x"fc",  x"eb",  x"21",  x"70",  x"33",  x"01",  x"31", -- 0038
         x"00",  x"ed",  x"b0",  x"eb",  x"01",  x"4f",  x"00",  x"09", -- 0040
         x"eb",  x"21",  x"a1",  x"33",  x"01",  x"33",  x"00",  x"ed", -- 0048
         x"b0",  x"eb",  x"01",  x"4d",  x"00",  x"09",  x"eb",  x"21", -- 0050
         x"d7",  x"33",  x"01",  x"39",  x"00",  x"ed",  x"b0",  x"eb", -- 0058
         x"01",  x"47",  x"00",  x"09",  x"eb",  x"21",  x"18",  x"34", -- 0060
         x"01",  x"22",  x"00",  x"ed",  x"b0",  x"eb",  x"01",  x"5e", -- 0068
         x"00",  x"09",  x"eb",  x"21",  x"3a",  x"34",  x"01",  x"10", -- 0070
         x"00",  x"ed",  x"b0",  x"eb",  x"01",  x"70",  x"00",  x"09", -- 0078
         x"eb",  x"21",  x"4b",  x"34",  x"01",  x"38",  x"00",  x"ed", -- 0080
         x"b0",  x"eb",  x"01",  x"54",  x"00",  x"09",  x"eb",  x"21", -- 0088
         x"0a",  x"03",  x"01",  x"1c",  x"00",  x"ed",  x"b0",  x"11", -- 0090
         x"92",  x"0c",  x"21",  x"5e",  x"33",  x"01",  x"12",  x"00", -- 0098
         x"ed",  x"b0",  x"3e",  x"01",  x"32",  x"c7",  x"0c",  x"cd", -- 00A0
         x"60",  x"2a",  x"3a",  x"03",  x"0c",  x"fe",  x"55",  x"28", -- 00A8
         x"08",  x"cd",  x"9a",  x"01",  x"c2",  x"f1",  x"00",  x"18", -- 00B0
         x"f1",  x"cd",  x"52",  x"33",  x"cd",  x"65",  x"32",  x"21", -- 00B8
         x"94",  x"3f",  x"cd",  x"e0",  x"01",  x"3e",  x"c0",  x"32", -- 00C0
         x"56",  x"0c",  x"2a",  x"00",  x"0c",  x"23",  x"22",  x"00", -- 00C8
         x"0c",  x"3e",  x"01",  x"32",  x"c7",  x"0c",  x"32",  x"c5", -- 00D0
         x"0c",  x"3e",  x"73",  x"32",  x"c8",  x"0c",  x"3e",  x"03", -- 00D8
         x"32",  x"1a",  x"0c",  x"3e",  x"14",  x"32",  x"e6",  x"0c", -- 00E0
         x"32",  x"e5",  x"0c",  x"32",  x"e4",  x"0c",  x"3a",  x"56", -- 00E8
         x"0c",  x"32",  x"bf",  x"0c",  x"cd",  x"e0",  x"29",  x"3a", -- 00F0
         x"e4",  x"0c",  x"b7",  x"ca",  x"79",  x"29",  x"3a",  x"c8", -- 00F8
         x"0c",  x"b7",  x"28",  x"42",  x"3e",  x"ff",  x"32",  x"56", -- 0100
         x"0c",  x"cd",  x"4a",  x"2a",  x"21",  x"80",  x"fb",  x"01", -- 0108
         x"bf",  x"00",  x"cd",  x"12",  x"32",  x"21",  x"3f",  x"3f", -- 0110
         x"cd",  x"d4",  x"01",  x"06",  x"05",  x"c5",  x"11",  x"d4", -- 0118
         x"fb",  x"21",  x"85",  x"34",  x"01",  x"14",  x"00",  x"ed", -- 0120
         x"b0",  x"0e",  x"c0",  x"cd",  x"ca",  x"01",  x"21",  x"d4", -- 0128
         x"fb",  x"01",  x"14",  x"00",  x"cd",  x"12",  x"32",  x"0e", -- 0130
         x"c0",  x"cd",  x"ca",  x"01",  x"c1",  x"10",  x"de",  x"af", -- 0138
         x"32",  x"03",  x"0c",  x"c3",  x"f1",  x"00",  x"3a",  x"56", -- 0140
         x"0c",  x"d6",  x"0a",  x"30",  x"02",  x"3e",  x"0a",  x"32", -- 0148
         x"56",  x"0c",  x"cd",  x"b2",  x"29",  x"21",  x"d1",  x"0c", -- 0150
         x"11",  x"d2",  x"0c",  x"af",  x"77",  x"01",  x"0e",  x"00", -- 0158
         x"ed",  x"b0",  x"21",  x"6f",  x"3f",  x"cd",  x"e0",  x"01", -- 0160
         x"cd",  x"97",  x"2e",  x"cd",  x"52",  x"33",  x"cd",  x"60", -- 0168
         x"2a",  x"3e",  x"73",  x"32",  x"c8",  x"0c",  x"c3",  x"f4", -- 0170
         x"28",  x"3a",  x"1a",  x"0c",  x"3d",  x"fe",  x"00",  x"28", -- 0178
         x"05",  x"fe",  x"04",  x"38",  x"07",  x"af",  x"32",  x"1a", -- 0180
         x"0c",  x"c3",  x"04",  x"29",  x"32",  x"1a",  x"0c",  x"cd", -- 0188
         x"65",  x"32",  x"21",  x"4e",  x"3f",  x"cd",  x"e0",  x"01", -- 0190
         x"3a",  x"1a",  x"0c",  x"b7",  x"ca",  x"04",  x"29",  x"3a", -- 0198
         x"e5",  x"0c",  x"32",  x"e6",  x"0c",  x"cb",  x"3f",  x"d6", -- 01A0
         x"03",  x"cd",  x"bb",  x"29",  x"cd",  x"65",  x"32",  x"c3", -- 01A8
         x"f4",  x"28",  x"3a",  x"e6",  x"0c",  x"32",  x"e5",  x"0c", -- 01B0
         x"3a",  x"e4",  x"0c",  x"4f",  x"3a",  x"e5",  x"0c",  x"fe", -- 01B8
         x"e0",  x"30",  x"07",  x"30",  x"0e",  x"3a",  x"e5",  x"0c", -- 01C0
         x"18",  x"09",  x"79",  x"c6",  x"05",  x"fe",  x"14",  x"38", -- 01C8
         x"02",  x"3e",  x"14",  x"32",  x"e4",  x"0c",  x"32",  x"e5", -- 01D0
         x"0c",  x"3a",  x"56",  x"0c",  x"32",  x"bf",  x"0c",  x"c9", -- 01D8
         x"cd",  x"56",  x"32",  x"3e",  x"d0",  x"cd",  x"ca",  x"01", -- 01E0
         x"21",  x"43",  x"0c",  x"36",  x"02",  x"cd",  x"65",  x"32", -- 01E8
         x"3a",  x"bf",  x"0c",  x"b7",  x"20",  x"10",  x"3a",  x"56", -- 01F0
         x"0c",  x"32",  x"bf",  x"0c",  x"3a",  x"e4",  x"0c",  x"3d", -- 01F8
         x"30",  x"01",  x"af",  x"32",  x"e4",  x"0c",  x"3a",  x"59", -- 0200
         x"0c",  x"b7",  x"20",  x"13",  x"af",  x"32",  x"cd",  x"0c", -- 0208
         x"21",  x"6d",  x"0c",  x"cb",  x"96",  x"21",  x"73",  x"0c", -- 0210
         x"cb",  x"96",  x"21",  x"79",  x"0c",  x"cb",  x"96",  x"cd", -- 0218
         x"c7",  x"01",  x"cd",  x"c7",  x"01",  x"cd",  x"97",  x"2b", -- 0220
         x"3a",  x"1a",  x"0c",  x"b7",  x"28",  x"1c",  x"3a",  x"c8", -- 0228
         x"0c",  x"b7",  x"c8",  x"3a",  x"e4",  x"0c",  x"b7",  x"c8", -- 0230
         x"21",  x"44",  x"0c",  x"af",  x"be",  x"28",  x"01",  x"35", -- 0238
         x"cd",  x"bb",  x"2e",  x"3a",  x"1a",  x"0c",  x"b7",  x"20", -- 0240
         x"a4",  x"c9",  x"2a",  x"18",  x"0c",  x"ed",  x"5b",  x"08", -- 0248
         x"0c",  x"b7",  x"ed",  x"52",  x"38",  x"06",  x"2a",  x"18", -- 0250
         x"0c",  x"22",  x"08",  x"0c",  x"cd",  x"56",  x"32",  x"c9", -- 0258
         x"21",  x"a8",  x"2a",  x"11",  x"68",  x"0c",  x"01",  x"12", -- 0260
         x"00",  x"ed",  x"b0",  x"3a",  x"c7",  x"0c",  x"47",  x"21", -- 0268
         x"68",  x"0c",  x"22",  x"93",  x"0c",  x"22",  x"97",  x"0c", -- 0270
         x"11",  x"00",  x"f8",  x"cd",  x"92",  x"0c",  x"19",  x"cd", -- 0278
         x"96",  x"0c",  x"2a",  x"93",  x"0c",  x"23",  x"23",  x"23", -- 0280
         x"23",  x"23",  x"23",  x"10",  x"e5",  x"cd",  x"ba",  x"2a", -- 0288
         x"c9",  x"22",  x"93",  x"0c",  x"22",  x"97",  x"0c",  x"11", -- 0290
         x"00",  x"f8",  x"cd",  x"92",  x"0c",  x"19",  x"cd",  x"96", -- 0298
         x"0c",  x"2a",  x"93",  x"0c",  x"cd",  x"30",  x"2b",  x"c9", -- 02A0
         x"da",  x"02",  x"1a",  x"0b",  x"00",  x"02",  x"dc",  x"02", -- 02A8
         x"1c",  x"0b",  x"00",  x"02",  x"de",  x"02",  x"1e",  x"0b", -- 02B0
         x"00",  x"02",  x"3a",  x"c7",  x"0c",  x"47",  x"21",  x"68", -- 02B8
         x"0c",  x"22",  x"93",  x"0c",  x"cd",  x"30",  x"2b",  x"2a", -- 02C0
         x"93",  x"0c",  x"c5",  x"cd",  x"a3",  x"32",  x"c1",  x"23", -- 02C8
         x"23",  x"23",  x"23",  x"23",  x"23",  x"10",  x"ea",  x"cd", -- 02D0
         x"de",  x"2a",  x"cd",  x"96",  x"32",  x"c9",  x"21",  x"c7", -- 02D8
         x"02",  x"11",  x"00",  x"f8",  x"19",  x"22",  x"c9",  x"0c", -- 02E0
         x"22",  x"cb",  x"0c",  x"3e",  x"1d",  x"32",  x"cf",  x"0c", -- 02E8
         x"3e",  x"17",  x"32",  x"ce",  x"0c",  x"af",  x"32",  x"e1", -- 02F0
         x"0c",  x"3a",  x"e1",  x"0c",  x"3c",  x"32",  x"e1",  x"0c", -- 02F8
         x"cb",  x"57",  x"20",  x"12",  x"2a",  x"cb",  x"0c",  x"36", -- 0300
         x"ea",  x"23",  x"36",  x"ec",  x"11",  x"3f",  x"00",  x"19", -- 0308
         x"36",  x"eb",  x"23",  x"36",  x"ed",  x"c9",  x"2a",  x"cb", -- 0310
         x"0c",  x"36",  x"ea",  x"cb",  x"5f",  x"28",  x"04",  x"af", -- 0318
         x"32",  x"e1",  x"0c",  x"23",  x"36",  x"ee",  x"11",  x"3f", -- 0320
         x"00",  x"19",  x"36",  x"eb",  x"23",  x"36",  x"ef",  x"c9", -- 0328
         x"2a",  x"93",  x"0c",  x"11",  x"05",  x"00",  x"19",  x"cb", -- 0330
         x"46",  x"28",  x"1c",  x"cb",  x"86",  x"cb",  x"4e",  x"20", -- 0338
         x"32",  x"cb",  x"56",  x"20",  x"2e",  x"cd",  x"92",  x"0c", -- 0340
         x"36",  x"f0",  x"23",  x"36",  x"f2",  x"11",  x"3f",  x"00", -- 0348
         x"19",  x"36",  x"f1",  x"23",  x"36",  x"f3",  x"c9",  x"cb", -- 0350
         x"c6",  x"cb",  x"4e",  x"20",  x"28",  x"cb",  x"56",  x"20", -- 0358
         x"24",  x"cd",  x"92",  x"0c",  x"36",  x"f4",  x"23",  x"36", -- 0360
         x"f6",  x"11",  x"3f",  x"00",  x"19",  x"36",  x"f5",  x"23", -- 0368
         x"36",  x"f7",  x"c9",  x"cd",  x"92",  x"0c",  x"36",  x"f8", -- 0370
         x"23",  x"36",  x"fe",  x"11",  x"3f",  x"00",  x"19",  x"36", -- 0378
         x"f9",  x"23",  x"36",  x"fb",  x"c9",  x"cd",  x"92",  x"0c", -- 0380
         x"36",  x"fc",  x"23",  x"36",  x"fe",  x"11",  x"3f",  x"00", -- 0388
         x"19",  x"36",  x"fd",  x"23",  x"36",  x"ff",  x"c9",  x"21", -- 0390
         x"1a",  x"0c",  x"af",  x"be",  x"20",  x"01",  x"c9",  x"3a", -- 0398
         x"cd",  x"0c",  x"cb",  x"bf",  x"32",  x"cd",  x"0c",  x"db", -- 03A0
         x"84",  x"ee",  x"00",  x"01",  x"40",  x"00",  x"2a",  x"cb", -- 03A8
         x"0c",  x"22",  x"c9",  x"0c",  x"32",  x"e2",  x"0c",  x"cb", -- 03B0
         x"4f",  x"ca",  x"6d",  x"2c",  x"3a",  x"e2",  x"0c",  x"2a", -- 03B8
         x"cb",  x"0c",  x"cb",  x"57",  x"ca",  x"d1",  x"2c",  x"3a", -- 03C0
         x"e2",  x"0c",  x"2a",  x"cb",  x"0c",  x"cb",  x"5f",  x"ca", -- 03C8
         x"37",  x"2d",  x"3a",  x"e2",  x"0c",  x"2a",  x"cb",  x"0c", -- 03D0
         x"cb",  x"67",  x"ca",  x"8c",  x"2d",  x"c3",  x"13",  x"2c", -- 03D8
         x"22",  x"cb",  x"0c",  x"2a",  x"c9",  x"0c",  x"cd",  x"28", -- 03E0
         x"32",  x"2a",  x"cb",  x"0c",  x"cd",  x"f9",  x"2a",  x"3a", -- 03E8
         x"cd",  x"0c",  x"cb",  x"7f",  x"3a",  x"c8",  x"0c",  x"b7", -- 03F0
         x"28",  x"04",  x"cd",  x"96",  x"32",  x"c9",  x"3a",  x"c5"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
