library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_8400 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_8400;

architecture rtl of rom1_8400 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"21",  x"52",  x"8c",  x"11",  x"4b",  x"fa",  x"3e",  x"2c", -- 0000
         x"cd",  x"24",  x"8a",  x"21",  x"5a",  x"8d",  x"11",  x"50", -- 0008
         x"fc",  x"01",  x"0e",  x"00",  x"ed",  x"b0",  x"06",  x"06", -- 0010
         x"21",  x"68",  x"8d",  x"11",  x"d0",  x"fc",  x"3e",  x"23", -- 0018
         x"cd",  x"24",  x"8a",  x"21",  x"18",  x"0c",  x"11",  x"19", -- 0020
         x"0c",  x"01",  x"90",  x"01",  x"36",  x"00",  x"ed",  x"b0", -- 0028
         x"11",  x"e8",  x"0c",  x"21",  x"38",  x"8b",  x"01",  x"12", -- 0030
         x"00",  x"ed",  x"b0",  x"3e",  x"02",  x"32",  x"1d",  x"0d", -- 0038
         x"3e",  x"02",  x"32",  x"1a",  x"0c",  x"cd",  x"73",  x"85", -- 0040
         x"3a",  x"03",  x"0c",  x"fe",  x"55",  x"28",  x"08",  x"cd", -- 0048
         x"9a",  x"01",  x"c2",  x"f1",  x"00",  x"18",  x"f1",  x"cd", -- 0050
         x"8f",  x"8b",  x"cd",  x"53",  x"8b",  x"21",  x"6e",  x"83", -- 0058
         x"cd",  x"e0",  x"01",  x"c5",  x"73",  x"85",  x"3e",  x"aa", -- 0060
         x"32",  x"56",  x"0c",  x"2a",  x"00",  x"0c",  x"23",  x"22", -- 0068
         x"00",  x"0c",  x"21",  x"00",  x"00",  x"af",  x"32",  x"42", -- 0070
         x"0d",  x"32",  x"1e",  x"0d",  x"22",  x"18",  x"0c",  x"22", -- 0078
         x"44",  x"0d",  x"3e",  x"fa",  x"32",  x"3a",  x"0d",  x"cd", -- 0080
         x"44",  x"85",  x"3a",  x"3a",  x"0d",  x"fe",  x"00",  x"28", -- 0088
         x"12",  x"3a",  x"1e",  x"0d",  x"fe",  x"5a",  x"38",  x"ef", -- 0090
         x"3a",  x"1a",  x"0c",  x"3d",  x"fe",  x"00",  x"28",  x"4c", -- 0098
         x"32",  x"1a",  x"0c",  x"3a",  x"56",  x"0c",  x"d6",  x"01", -- 00A0
         x"30",  x"02",  x"3e",  x"0c",  x"32",  x"56",  x"0c",  x"3a", -- 00A8
         x"3a",  x"0d",  x"fe",  x"00",  x"20",  x"0a",  x"3e",  x"fa", -- 00B0
         x"32",  x"3a",  x"0d",  x"cd",  x"5a",  x"85",  x"18",  x"ca", -- 00B8
         x"3a",  x"1d",  x"0d",  x"fe",  x"02",  x"30",  x"05",  x"c6", -- 00C0
         x"01",  x"32",  x"1d",  x"0d",  x"21",  x"ba",  x"83",  x"cd", -- 00C8
         x"e0",  x"01",  x"af",  x"32",  x"42",  x"0d",  x"32",  x"1e", -- 00D0
         x"0d",  x"3a",  x"56",  x"0c",  x"c6",  x"1e",  x"32",  x"56", -- 00D8
         x"0c",  x"cd",  x"8f",  x"8b",  x"cd",  x"53",  x"8b",  x"cd", -- 00E0
         x"73",  x"85",  x"18",  x"96",  x"2a",  x"18",  x"0c",  x"ed", -- 00E8
         x"5b",  x"04",  x"0c",  x"b7",  x"ed",  x"52",  x"38",  x"06", -- 00F0
         x"2a",  x"18",  x"0c",  x"22",  x"04",  x"0c",  x"af",  x"32", -- 00F8
         x"1a",  x"0c",  x"cd",  x"f0",  x"89",  x"21",  x"ca",  x"fb", -- 0100
         x"01",  x"28",  x"00",  x"cd",  x"4a",  x"8b",  x"21",  x"84", -- 0108
         x"83",  x"cd",  x"d4",  x"01",  x"3e",  x"96",  x"32",  x"56", -- 0110
         x"0c",  x"06",  x"05",  x"c5",  x"11",  x"d8",  x"fb",  x"21", -- 0118
         x"3a",  x"8e",  x"01",  x"14",  x"00",  x"ed",  x"b0",  x"0e", -- 0120
         x"fa",  x"cd",  x"ca",  x"01",  x"21",  x"d8",  x"fb",  x"01", -- 0128
         x"14",  x"00",  x"cd",  x"4a",  x"8b",  x"0e",  x"fa",  x"cd", -- 0130
         x"ca",  x"01",  x"c1",  x"10",  x"de",  x"af",  x"32",  x"03", -- 0138
         x"0c",  x"c3",  x"f1",  x"00",  x"cd",  x"f0",  x"89",  x"3e", -- 0140
         x"c8",  x"cd",  x"ca",  x"01",  x"21",  x"43",  x"0c",  x"36", -- 0148
         x"02",  x"cd",  x"c7",  x"01",  x"cd",  x"c7",  x"01",  x"cd", -- 0150
         x"f0",  x"89",  x"cd",  x"51",  x"87",  x"cd",  x"76",  x"88", -- 0158
         x"3a",  x"1e",  x"0d",  x"fe",  x"5a",  x"d0",  x"3a",  x"3a", -- 0160
         x"0d",  x"d6",  x"02",  x"32",  x"3a",  x"0d",  x"fe",  x"00", -- 0168
         x"c8",  x"18",  x"de",  x"21",  x"a3",  x"85",  x"11",  x"68", -- 0170
         x"0c",  x"01",  x"0f",  x"00",  x"ed",  x"b0",  x"3a",  x"1d", -- 0178
         x"0d",  x"47",  x"21",  x"68",  x"0c",  x"22",  x"e9",  x"0c", -- 0180
         x"22",  x"ed",  x"0c",  x"11",  x"00",  x"f8",  x"cd",  x"e8", -- 0188
         x"0c",  x"19",  x"cd",  x"ec",  x"0c",  x"2a",  x"e9",  x"0c", -- 0190
         x"23",  x"23",  x"23",  x"23",  x"23",  x"10",  x"e6",  x"cd", -- 0198
         x"b2",  x"85",  x"c9",  x"88",  x"01",  x"09",  x"06",  x"00", -- 01A0
         x"90",  x"01",  x"11",  x"06",  x"00",  x"98",  x"01",  x"19", -- 01A8
         x"06",  x"00",  x"3a",  x"1d",  x"0d",  x"47",  x"21",  x"68", -- 01B0
         x"0c",  x"22",  x"e9",  x"0c",  x"cd",  x"40",  x"87",  x"2a", -- 01B8
         x"e9",  x"0c",  x"c5",  x"cd",  x"aa",  x"8b",  x"c1",  x"23", -- 01C0
         x"23",  x"23",  x"23",  x"23",  x"10",  x"eb",  x"cd",  x"d5", -- 01C8
         x"85",  x"cd",  x"9d",  x"8b",  x"c9",  x"21",  x"50",  x"07", -- 01D0
         x"11",  x"00",  x"f8",  x"19",  x"22",  x"1f",  x"0d",  x"22", -- 01D8
         x"21",  x"0d",  x"3e",  x"1d",  x"32",  x"25",  x"0d",  x"3a", -- 01E0
         x"0f",  x"00",  x"32",  x"24",  x"0d",  x"af",  x"32",  x"37", -- 01E8
         x"0d",  x"3a",  x"37",  x"0d",  x"3c",  x"32",  x"37",  x"0d", -- 01F0
         x"fe",  x"06",  x"30",  x"2a",  x"2a",  x"21",  x"0d",  x"cd", -- 01F8
         x"51",  x"86",  x"3a",  x"25",  x"0d",  x"fe",  x"1d",  x"38", -- 0200
         x"06",  x"3a",  x"1e",  x"0d",  x"fe",  x"24",  x"d0",  x"3a", -- 0208
         x"3d",  x"0d",  x"cb",  x"4f",  x"28",  x"09",  x"36",  x"d5", -- 0210
         x"2b",  x"36",  x"d4",  x"cd",  x"71",  x"89",  x"c9",  x"36", -- 0218
         x"d3",  x"2b",  x"36",  x"d2",  x"18",  x"f5",  x"2a",  x"21", -- 0220
         x"0d",  x"fe",  x"0c",  x"38",  x"04",  x"af",  x"32",  x"37", -- 0228
         x"0d",  x"cd",  x"51",  x"86",  x"3a",  x"25",  x"0d",  x"fe", -- 0230
         x"1d",  x"38",  x"06",  x"3a",  x"1e",  x"0d",  x"fe",  x"24", -- 0238
         x"d0",  x"36",  x"dc",  x"2b",  x"3a",  x"3d",  x"0d",  x"cb", -- 0240
         x"4f",  x"28",  x"02",  x"18",  x"cc",  x"36",  x"d2",  x"18", -- 0248
         x"ca",  x"3a",  x"25",  x"0d",  x"fe",  x"1d",  x"38",  x"0a", -- 0250
         x"3a",  x"1e",  x"0d",  x"fe",  x"48",  x"38",  x"03",  x"2b", -- 0258
         x"18",  x"18",  x"36",  x"d1",  x"2b",  x"3a",  x"43",  x"0d", -- 0260
         x"cb",  x"47",  x"28",  x"0e",  x"36",  x"00",  x"cd",  x"cf", -- 0268
         x"8a",  x"36",  x"00",  x"cb",  x"87",  x"32",  x"43",  x"0d", -- 0270
         x"18",  x"03",  x"cd",  x"cf",  x"8a",  x"23",  x"36",  x"d0", -- 0278
         x"23",  x"3a",  x"42",  x"0d",  x"fe",  x"01",  x"38",  x"16", -- 0280
         x"fe",  x"03",  x"38",  x"1b",  x"fe",  x"05",  x"38",  x"20", -- 0288
         x"fe",  x"08",  x"38",  x"25",  x"fe",  x"0c",  x"38",  x"25", -- 0290
         x"fe",  x"0e",  x"38",  x"25",  x"18",  x"27",  x"cd",  x"ce", -- 0298
         x"86",  x"3e",  x"d7",  x"cd",  x"da",  x"86",  x"c9",  x"cd", -- 02A0
         x"ce",  x"86",  x"3e",  x"d9",  x"cd",  x"da",  x"86",  x"c9", -- 02A8
         x"cd",  x"ce",  x"86",  x"3e",  x"db",  x"cd",  x"da",  x"86", -- 02B0
         x"c9",  x"3e",  x"e2",  x"18",  x"0a",  x"3e",  x"e4",  x"18", -- 02B8
         x"06",  x"3e",  x"e6",  x"18",  x"02",  x"3e",  x"e8",  x"cd", -- 02C0
         x"d0",  x"86",  x"cd",  x"d8",  x"86",  x"c9",  x"3e",  x"e0", -- 02C8
         x"77",  x"23",  x"3c",  x"77",  x"cd",  x"cb",  x"8a",  x"c9", -- 02D0
         x"3e",  x"db",  x"4f",  x"3a",  x"25",  x"0d",  x"fe",  x"1d", -- 02D8
         x"38",  x"0a",  x"3a",  x"1e",  x"0d",  x"fe",  x"48",  x"38", -- 02E0
         x"03",  x"2b",  x"18",  x"05",  x"79",  x"77",  x"3d",  x"2b", -- 02E8
         x"77",  x"cd",  x"cb",  x"8a",  x"c9",  x"cd",  x"cf",  x"8a", -- 02F0
         x"2b",  x"36",  x"ee",  x"23",  x"36",  x"de",  x"23",  x"36", -- 02F8
         x"df",  x"23",  x"36",  x"00",  x"3a",  x"43",  x"0d",  x"cb", -- 0300
         x"c7",  x"32",  x"43",  x"0d",  x"3a",  x"25",  x"0d",  x"fe", -- 0308
         x"1d",  x"38",  x"06",  x"3a",  x"1e",  x"0d",  x"fe",  x"48", -- 0310
         x"d0",  x"cd",  x"cb",  x"8a",  x"36",  x"00",  x"2b",  x"36", -- 0318
         x"f4",  x"2b",  x"36",  x"f3",  x"2b",  x"36",  x"dd",  x"3a", -- 0320
         x"25",  x"0d",  x"fe",  x"1d",  x"38",  x"06",  x"3a",  x"1e", -- 0328
         x"0d",  x"fe",  x"24",  x"d0",  x"cd",  x"cb",  x"8a",  x"23", -- 0330
         x"36",  x"d4",  x"23",  x"36",  x"d5",  x"c3",  x"1b",  x"86", -- 0338
         x"2a",  x"e9",  x"0c",  x"11",  x"04",  x"00",  x"19",  x"3e", -- 0340
         x"ff",  x"be",  x"c8",  x"cd",  x"e8",  x"0c",  x"36",  x"ef", -- 0348
         x"c9",  x"21",  x"43",  x"0c",  x"35",  x"c0",  x"36",  x"02", -- 0350
         x"3a",  x"1d",  x"0d",  x"47",  x"21",  x"68",  x"0c",  x"22", -- 0358
         x"e9",  x"0c",  x"22",  x"ed",  x"0c",  x"c5",  x"cd",  x"7e", -- 0360
         x"87",  x"c1",  x"2a",  x"e9",  x"0c",  x"3a",  x"1e",  x"0d", -- 0368
         x"fe",  x"5a",  x"d0",  x"23",  x"23",  x"23",  x"23",  x"23", -- 0370
         x"10",  x"e5",  x"cd",  x"89",  x"89",  x"c9",  x"2a",  x"e9", -- 0378
         x"0c",  x"23",  x"23",  x"23",  x"23",  x"db",  x"83",  x"32", -- 0380
         x"26",  x"0d",  x"7e",  x"fe",  x"00",  x"20",  x"09",  x"3a", -- 0388
         x"26",  x"0d",  x"fe",  x"5a",  x"38",  x"02",  x"36",  x"01", -- 0390
         x"7e",  x"2b",  x"2b",  x"2b",  x"2b",  x"fe",  x"01",  x"20", -- 0398
         x"04",  x"cd",  x"b7",  x"87",  x"c8",  x"cd",  x"e8",  x"0c", -- 03A0
         x"36",  x"00",  x"cd",  x"d4",  x"8b",  x"cd",  x"e8",  x"0c", -- 03A8
         x"cd",  x"40",  x"87",  x"cd",  x"71",  x"89",  x"c9",  x"cd", -- 03B0
         x"c6",  x"87",  x"c8",  x"2a",  x"e9",  x"0c",  x"23",  x"23", -- 03B8
         x"23",  x"34",  x"2b",  x"2b",  x"2b",  x"c9",  x"cd",  x"e8", -- 03C0
         x"0c",  x"cd",  x"cb",  x"8a",  x"7e",  x"e6",  x"f0",  x"fe", -- 03C8
         x"e0",  x"28",  x"39",  x"fe",  x"c0",  x"d8",  x"3a",  x"1e", -- 03D0
         x"0d",  x"3c",  x"32",  x"1e",  x"0d",  x"21",  x"98",  x"83", -- 03D8
         x"cd",  x"d4",  x"01",  x"cd",  x"f0",  x"89",  x"cd",  x"e8", -- 03E0
         x"0c",  x"36",  x"00",  x"2a",  x"e9",  x"0c",  x"23",  x"23", -- 03E8
         x"3a",  x"26",  x"0d",  x"e6",  x"37",  x"fe",  x"12",  x"30", -- 03F0
         x"02",  x"c6",  x"0c",  x"77",  x"23",  x"36",  x"06",  x"23"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
