library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_8800 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_8800;

architecture rtl of rom1_8800 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"36",  x"00",  x"cd",  x"d4",  x"8b",  x"cd",  x"40",  x"87", -- 0000
         x"3e",  x"01",  x"3d",  x"c9",  x"2a",  x"18",  x"0c",  x"3a", -- 0008
         x"42",  x"0d",  x"fe",  x"0f",  x"38",  x"11",  x"21",  x"ac", -- 0010
         x"83",  x"cd",  x"d4",  x"01",  x"f5",  x"3a",  x"1e",  x"0d", -- 0018
         x"3c",  x"32",  x"1e",  x"0d",  x"f1",  x"18",  x"bc",  x"11", -- 0020
         x"05",  x"00",  x"19",  x"22",  x"18",  x"0c",  x"2a",  x"44", -- 0028
         x"0d",  x"19",  x"22",  x"44",  x"0d",  x"3c",  x"32",  x"42", -- 0030
         x"0d",  x"cd",  x"f0",  x"89",  x"21",  x"91",  x"83",  x"cd", -- 0038
         x"d4",  x"01",  x"cd",  x"47",  x"88",  x"18",  x"9c",  x"2a", -- 0040
         x"44",  x"0d",  x"11",  x"dc",  x"05",  x"b7",  x"ed",  x"52", -- 0048
         x"d8",  x"21",  x"00",  x"00",  x"22",  x"44",  x"0d",  x"3a", -- 0050
         x"1a",  x"0c",  x"fe",  x"04",  x"d0",  x"3c",  x"32",  x"1a", -- 0058
         x"0c",  x"cd",  x"f0",  x"89",  x"21",  x"b1",  x"83",  x"cd", -- 0060
         x"e0",  x"01",  x"c9",  x"21",  x"84",  x"fb",  x"3e",  x"f0", -- 0068
         x"06",  x"06",  x"cd",  x"9d",  x"8a",  x"c9",  x"cd",  x"6b", -- 0070
         x"88",  x"2a",  x"21",  x"0d",  x"22",  x"1f",  x"0d",  x"db", -- 0078
         x"84",  x"ee",  x"00",  x"32",  x"3d",  x"0d",  x"cb",  x"47", -- 0080
         x"ca",  x"05",  x"89",  x"cb",  x"67",  x"cc",  x"d8",  x"88", -- 0088
         x"cb",  x"5f",  x"cc",  x"cb",  x"88",  x"cb",  x"57",  x"ca", -- 0090
         x"bc",  x"88",  x"cb",  x"4f",  x"cc",  x"a3",  x"88",  x"cd", -- 0098
         x"e9",  x"88",  x"c9",  x"e5",  x"06",  x"02",  x"cd",  x"bd", -- 00A0
         x"8a",  x"23",  x"7e",  x"e1",  x"fe",  x"f2",  x"20",  x"36", -- 00A8
         x"23",  x"23",  x"23",  x"7e",  x"2b",  x"2b",  x"fe",  x"ed", -- 00B0
         x"20",  x"2c",  x"18",  x"2d",  x"2b",  x"7e",  x"fe",  x"f0", -- 00B8
         x"28",  x"27",  x"2b",  x"7e",  x"23",  x"fe",  x"f2",  x"20", -- 00C0
         x"1d",  x"18",  x"1e",  x"2b",  x"2b",  x"7e",  x"23",  x"fe", -- 00C8
         x"f2",  x"20",  x"16",  x"cd",  x"cf",  x"8a",  x"18",  x"0e", -- 00D0
         x"06",  x"02",  x"cd",  x"bd",  x"8a",  x"23",  x"7e",  x"cd", -- 00D8
         x"cf",  x"8a",  x"fe",  x"f2",  x"28",  x"03",  x"22",  x"21", -- 00E0
         x"0d",  x"2a",  x"1f",  x"0d",  x"cd",  x"d3",  x"8a",  x"2a", -- 00E8
         x"21",  x"0d",  x"22",  x"1f",  x"0d",  x"cd",  x"f1",  x"85", -- 00F0
         x"cd",  x"9d",  x"8b",  x"cd",  x"6b",  x"88",  x"3a",  x"3d", -- 00F8
         x"0d",  x"2a",  x"21",  x"0d",  x"c9",  x"cd",  x"9d",  x"8b", -- 0100
         x"cd",  x"f5",  x"86",  x"3a",  x"24",  x"0d",  x"fe",  x"07", -- 0108
         x"38",  x"33",  x"2a",  x"18",  x"0c",  x"3a",  x"42",  x"0d", -- 0110
         x"fe",  x"00",  x"c8",  x"5f",  x"16",  x"00",  x"b7",  x"ed", -- 0118
         x"52",  x"30",  x"03",  x"21",  x"00",  x"00",  x"22",  x"18", -- 0120
         x"0c",  x"3a",  x"42",  x"0d",  x"5f",  x"3a",  x"1e",  x"0d", -- 0128
         x"83",  x"32",  x"1e",  x"0d",  x"cd",  x"f0",  x"89",  x"cd", -- 0130
         x"89",  x"89",  x"21",  x"9f",  x"83",  x"cd",  x"d4",  x"01", -- 0138
         x"af",  x"32",  x"42",  x"0d",  x"c9",  x"2a",  x"18",  x"0c", -- 0140
         x"3a",  x"42",  x"0d",  x"fe",  x"00",  x"c8",  x"5f",  x"16", -- 0148
         x"00",  x"19",  x"19",  x"19",  x"22",  x"18",  x"0c",  x"2a", -- 0150
         x"44",  x"0d",  x"19",  x"19",  x"19",  x"22",  x"44",  x"0d", -- 0158
         x"af",  x"32",  x"42",  x"0d",  x"cd",  x"f0",  x"89",  x"21", -- 0160
         x"b1",  x"83",  x"cd",  x"d4",  x"01",  x"cd",  x"47",  x"88", -- 0168
         x"c9",  x"3a",  x"1e",  x"0d",  x"21",  x"8f",  x"ff",  x"06", -- 0170
         x"2c",  x"fe",  x"24",  x"d4",  x"c5",  x"89",  x"21",  x"4e", -- 0178
         x"ff",  x"06",  x"2d",  x"fe",  x"48",  x"d4",  x"c5",  x"89", -- 0180
         x"c9",  x"cd",  x"71",  x"89",  x"fe",  x"24",  x"38",  x"15", -- 0188
         x"fe",  x"48",  x"38",  x"1a",  x"fe",  x"62",  x"38",  x"02", -- 0190
         x"3e",  x"61",  x"d6",  x"48",  x"21",  x"0d",  x"ff",  x"06", -- 0198
         x"2e",  x"cd",  x"b9",  x"89",  x"c9",  x"21",  x"8f",  x"ff", -- 01A0
         x"06",  x"2c",  x"cd",  x"b9",  x"89",  x"c9",  x"21",  x"4e", -- 01A8
         x"ff",  x"d6",  x"24",  x"06",  x"2d",  x"cd",  x"b9",  x"89", -- 01B0
         x"c9",  x"0e",  x"c7",  x"fe",  x"04",  x"d8",  x"d6",  x"04", -- 01B8
         x"38",  x"05",  x"0c",  x"18",  x"f9",  x"0e",  x"cf",  x"71", -- 01C0
         x"23",  x"10",  x"fc",  x"c9",  x"21",  x"f5",  x"8b",  x"11", -- 01C8
         x"00",  x"f8",  x"01",  x"40",  x"00",  x"ed",  x"b0",  x"21", -- 01D0
         x"05",  x"f9",  x"3e",  x"eb",  x"06",  x"35",  x"cd",  x"93", -- 01D8
         x"8a",  x"21",  x"0b",  x"f8",  x"22",  x"3f",  x"0c",  x"2a", -- 01E0
         x"04",  x"0c",  x"22",  x"3d",  x"0c",  x"cd",  x"70",  x"02", -- 01E8
         x"21",  x"1b",  x"f8",  x"22",  x"3f",  x"0c",  x"2a",  x"18", -- 01F0
         x"0c",  x"22",  x"3d",  x"0c",  x"cd",  x"70",  x"02",  x"21", -- 01F8
         x"2a",  x"f8",  x"22",  x"3f",  x"0c",  x"3a",  x"1a",  x"0c", -- 0200
         x"6f",  x"26",  x"00",  x"22",  x"3d",  x"0c",  x"cd",  x"70", -- 0208
         x"02",  x"21",  x"3b",  x"f8",  x"22",  x"3f",  x"0c",  x"26", -- 0210
         x"00",  x"3a",  x"1e",  x"0d",  x"6f",  x"22",  x"3d",  x"0c", -- 0218
         x"cd",  x"70",  x"02",  x"c9",  x"c5",  x"d5",  x"e5",  x"06", -- 0220
         x"00",  x"4f",  x"ed",  x"b0",  x"e1",  x"5f",  x"16",  x"00", -- 0228
         x"19",  x"d1",  x"eb",  x"01",  x"40",  x"00",  x"09",  x"eb", -- 0230
         x"c1",  x"10",  x"e9",  x"c9",  x"21",  x"3c",  x"f8",  x"3e", -- 0238
         x"f2",  x"06",  x"1f",  x"cd",  x"9d",  x"8a",  x"06",  x"38", -- 0240
         x"cd",  x"98",  x"8a",  x"06",  x"0c",  x"cd",  x"a5",  x"8a", -- 0248
         x"06",  x"06",  x"3e",  x"f0",  x"cd",  x"a5",  x"8a",  x"3e", -- 0250
         x"f2",  x"21",  x"04",  x"f8",  x"06",  x"0e",  x"cd",  x"9d", -- 0258
         x"8a",  x"21",  x"40",  x"fd",  x"3e",  x"f1",  x"06",  x"04", -- 0260
         x"cd",  x"93",  x"8a",  x"06",  x"39",  x"cd",  x"b8",  x"8a", -- 0268
         x"06",  x"03",  x"cd",  x"93",  x"8a",  x"21",  x"45",  x"fd", -- 0270
         x"cd",  x"23",  x"8b",  x"c9",  x"3e",  x"ea",  x"77",  x"06", -- 0278
         x"01",  x"cd",  x"bd",  x"8a",  x"77",  x"2b",  x"77",  x"06", -- 0280
         x"01",  x"cd",  x"bd",  x"8a",  x"2b",  x"77",  x"23",  x"77", -- 0288
         x"23",  x"77",  x"c9",  x"77",  x"23",  x"10",  x"fc",  x"c9", -- 0290
         x"77",  x"2b",  x"10",  x"fc",  x"c9",  x"77",  x"11",  x"40", -- 0298
         x"00",  x"19",  x"10",  x"f9",  x"c9",  x"77",  x"11",  x"40", -- 02A0
         x"00",  x"b7",  x"ed",  x"52",  x"10",  x"f7",  x"c9",  x"11", -- 02A8
         x"40",  x"00",  x"b7",  x"ed",  x"52",  x"10",  x"f8",  x"c9", -- 02B0
         x"48",  x"06",  x"00",  x"09",  x"c9",  x"11",  x"40",  x"00", -- 02B8
         x"19",  x"10",  x"fa",  x"c9",  x"48",  x"06",  x"00",  x"b7", -- 02C0
         x"ed",  x"42",  x"c9",  x"06",  x"01",  x"18",  x"ee",  x"06", -- 02C8
         x"01",  x"18",  x"dc",  x"e5",  x"cd",  x"cf",  x"8a",  x"af", -- 02D0
         x"06",  x"03",  x"cd",  x"93",  x"8a",  x"cd",  x"cb",  x"8a", -- 02D8
         x"2b",  x"3a",  x"25",  x"0d",  x"fe",  x"1d",  x"38",  x"07", -- 02E0
         x"3a",  x"1e",  x"0d",  x"fe",  x"48",  x"30",  x"1e",  x"af", -- 02E8
         x"06",  x"03",  x"cd",  x"98",  x"8a",  x"23",  x"cd",  x"cb", -- 02F0
         x"8a",  x"3a",  x"25",  x"0d",  x"fe",  x"1d",  x"38",  x"07", -- 02F8
         x"3a",  x"1e",  x"0d",  x"fe",  x"24",  x"30",  x"06",  x"af", -- 0300
         x"06",  x"02",  x"cd",  x"93",  x"8a",  x"e1",  x"3a",  x"43", -- 0308
         x"0d",  x"cb",  x"47",  x"c8",  x"cb",  x"87",  x"32",  x"43", -- 0310
         x"0d",  x"e5",  x"af",  x"2b",  x"77",  x"cd",  x"cf",  x"8a", -- 0318
         x"77",  x"e1",  x"c9",  x"3e",  x"f2",  x"06",  x"01",  x"0e", -- 0320
         x"0a",  x"c5",  x"e5",  x"cd",  x"93",  x"8a",  x"e1",  x"cd", -- 0328
         x"cb",  x"8a",  x"c1",  x"04",  x"0d",  x"20",  x"f2",  x"c9", -- 0330
         x"2a",  x"00",  x"00",  x"c9",  x"22",  x"00",  x"00",  x"c9", -- 0338
         x"ed",  x"5b",  x"00",  x"00",  x"c9",  x"ed",  x"53",  x"00", -- 0340
         x"00",  x"c9",  x"54",  x"5d",  x"13",  x"36",  x"00",  x"0b", -- 0348
         x"ed",  x"b0",  x"c9",  x"cd",  x"3c",  x"8a",  x"cd",  x"cc", -- 0350
         x"89",  x"21",  x"7c",  x"f9",  x"06",  x"38",  x"3e",  x"f2", -- 0358
         x"cd",  x"98",  x"8a",  x"21",  x"7b",  x"f8",  x"3e",  x"ed", -- 0360
         x"06",  x"01",  x"cd",  x"9d",  x"8a",  x"3e",  x"ec",  x"06", -- 0368
         x"02",  x"cd",  x"9d",  x"8a",  x"3e",  x"ed",  x"06",  x"1c", -- 0370
         x"cd",  x"9d",  x"8a",  x"21",  x"ba",  x"f8",  x"cd",  x"7c", -- 0378
         x"8a",  x"21",  x"40",  x"f8",  x"11",  x"41",  x"f8",  x"01", -- 0380
         x"3f",  x"00",  x"36",  x"00",  x"ed",  x"b0",  x"c9",  x"21", -- 0388
         x"00",  x"f8",  x"11",  x"01",  x"f8",  x"36",  x"00",  x"01", -- 0390
         x"ff",  x"07",  x"ed",  x"b0",  x"c9",  x"e5",  x"2a",  x"21", -- 0398
         x"0d",  x"cd",  x"bc",  x"8b",  x"ed",  x"43",  x"24",  x"0d", -- 03A0
         x"e1",  x"c9",  x"e5",  x"5e",  x"23",  x"56",  x"eb",  x"cd", -- 03A8
         x"bc",  x"8b",  x"e1",  x"23",  x"23",  x"71",  x"23",  x"70", -- 03B0
         x"2b",  x"2b",  x"2b",  x"c9",  x"11",  x"00",  x"f8",  x"01", -- 03B8
         x"00",  x"00",  x"b7",  x"ed",  x"52",  x"11",  x"40",  x"00", -- 03C0
         x"b7",  x"ed",  x"52",  x"c8",  x"38",  x"03",  x"04",  x"18", -- 03C8
         x"f7",  x"19",  x"4d",  x"c9",  x"2a",  x"e9",  x"0c",  x"23", -- 03D0
         x"23",  x"4e",  x"23",  x"46",  x"21",  x"00",  x"f8",  x"11", -- 03D8
         x"40",  x"00",  x"af",  x"b8",  x"28",  x"05",  x"05",  x"19", -- 03E0
         x"d8",  x"18",  x"f7",  x"09",  x"2b",  x"eb",  x"2a",  x"e9", -- 03E8
         x"0c",  x"73",  x"23",  x"72",  x"c9",  x"3d",  x"3d",  x"20", -- 03F0
         x"52",  x"45",  x"4b",  x"4f",  x"52",  x"44",  x"3a",  x"20"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
