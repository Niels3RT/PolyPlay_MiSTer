library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_5000 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_5000;

architecture rtl of rom1_5000 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"cd",  x"b7",  x"02",  x"cd",  x"55",  x"59",  x"cd",  x"ea", -- 0000
         x"59",  x"11",  x"00",  x"ec",  x"21",  x"6f",  x"5c",  x"3a", -- 0008
         x"db",  x"5f",  x"47",  x"c5",  x"4e",  x"23",  x"46",  x"23", -- 0010
         x"7e",  x"23",  x"eb",  x"09",  x"eb",  x"47",  x"c5",  x"01", -- 0018
         x"08",  x"00",  x"ed",  x"b0",  x"cd",  x"64",  x"59",  x"c1", -- 0020
         x"10",  x"f4",  x"e5",  x"d5",  x"eb",  x"01",  x"08",  x"00", -- 0028
         x"09",  x"eb",  x"21",  x"12",  x"0d",  x"cd",  x"64",  x"59", -- 0030
         x"d1",  x"e1",  x"c1",  x"10",  x"d6",  x"fd",  x"21",  x"01", -- 0038
         x"0d",  x"fd",  x"36",  x"00",  x"00",  x"3e",  x"02",  x"32", -- 0040
         x"00",  x"0d",  x"3e",  x"ff",  x"32",  x"56",  x"0c",  x"3e", -- 0048
         x"4d",  x"32",  x"bf",  x"0c",  x"3e",  x"07",  x"32",  x"46", -- 0050
         x"0d",  x"af",  x"32",  x"33",  x"0d",  x"32",  x"4a",  x"0d", -- 0058
         x"32",  x"49",  x"0d",  x"3e",  x"0f",  x"32",  x"32",  x"0d", -- 0060
         x"3e",  x"01",  x"32",  x"34",  x"0d",  x"3e",  x"20",  x"32", -- 0068
         x"3b",  x"0d",  x"3e",  x"c0",  x"32",  x"35",  x"0d",  x"21", -- 0070
         x"60",  x"ff",  x"22",  x"39",  x"0d",  x"21",  x"40",  x"00", -- 0078
         x"22",  x"3c",  x"0d",  x"3e",  x"01",  x"32",  x"3f",  x"0d", -- 0080
         x"3e",  x"03",  x"32",  x"40",  x"0d",  x"3e",  x"05",  x"32", -- 0088
         x"41",  x"0d",  x"3e",  x"08",  x"32",  x"42",  x"0d",  x"3e", -- 0090
         x"c6",  x"32",  x"43",  x"0d",  x"dd",  x"21",  x"37",  x"5c", -- 0098
         x"21",  x"00",  x"f8",  x"36",  x"20",  x"11",  x"01",  x"f8", -- 00A0
         x"01",  x"ff",  x"07",  x"ed",  x"b0",  x"cd",  x"0b",  x"57", -- 00A8
         x"17",  x"5a",  x"21",  x"0a",  x"f8",  x"22",  x"3f",  x"0c", -- 00B0
         x"2a",  x"0c",  x"0c",  x"22",  x"3d",  x"0c",  x"cd",  x"70", -- 00B8
         x"02",  x"21",  x"1a",  x"f8",  x"22",  x"3f",  x"0c",  x"2a", -- 00C0
         x"18",  x"0c",  x"22",  x"3d",  x"0c",  x"cd",  x"70",  x"02", -- 00C8
         x"fd",  x"cb",  x"00",  x"46",  x"28",  x"0a",  x"06",  x"40", -- 00D0
         x"21",  x"80",  x"ff",  x"36",  x"10",  x"23",  x"10",  x"fb", -- 00D8
         x"21",  x"01",  x"f9",  x"e5",  x"06",  x"04",  x"11",  x"40", -- 00E0
         x"00",  x"19",  x"36",  x"d0",  x"10",  x"fb",  x"e1",  x"06", -- 00E8
         x"14",  x"36",  x"d0",  x"23",  x"10",  x"fb",  x"2b",  x"06", -- 00F0
         x"04",  x"19",  x"36",  x"d0",  x"10",  x"fb",  x"06",  x"14", -- 00F8
         x"36",  x"d0",  x"2b",  x"10",  x"fb",  x"cd",  x"0b",  x"57", -- 0100
         x"59",  x"5a",  x"21",  x"57",  x"f9",  x"06",  x"10",  x"36", -- 0108
         x"10",  x"23",  x"10",  x"fb",  x"21",  x"d7",  x"f9",  x"06", -- 0110
         x"29",  x"36",  x"c8",  x"23",  x"10",  x"fb",  x"21",  x"17", -- 0118
         x"fa",  x"06",  x"29",  x"36",  x"c8",  x"23",  x"10",  x"fb", -- 0120
         x"21",  x"6b",  x"f9",  x"3a",  x"41",  x"0d",  x"06",  x"d8", -- 0128
         x"70",  x"23",  x"70",  x"cd",  x"2a",  x"57",  x"21",  x"7e", -- 0130
         x"fb",  x"70",  x"23",  x"70",  x"cd",  x"2a",  x"57",  x"21", -- 0138
         x"71",  x"f9",  x"3a",  x"40",  x"0d",  x"06",  x"d6",  x"70", -- 0140
         x"23",  x"70",  x"cd",  x"2a",  x"57",  x"fd",  x"cb",  x"00", -- 0148
         x"46",  x"28",  x"09",  x"21",  x"3e",  x"fc",  x"70",  x"23", -- 0150
         x"70",  x"cd",  x"2a",  x"57",  x"21",  x"77",  x"f9",  x"3a", -- 0158
         x"3f",  x"0d",  x"06",  x"da",  x"70",  x"23",  x"70",  x"cd", -- 0160
         x"2a",  x"57",  x"fd",  x"cb",  x"00",  x"46",  x"28",  x"18", -- 0168
         x"21",  x"fe",  x"fc",  x"70",  x"23",  x"70",  x"cd",  x"2a", -- 0170
         x"57",  x"2a",  x"39",  x"0d",  x"36",  x"c2",  x"23",  x"36", -- 0178
         x"c4",  x"01",  x"c0",  x"ff",  x"09",  x"22",  x"37",  x"0d", -- 0180
         x"21",  x"02",  x"0d",  x"3e",  x"20",  x"77",  x"54",  x"5d", -- 0188
         x"13",  x"01",  x"2f",  x"00",  x"ed",  x"b0",  x"11",  x"47", -- 0190
         x"5b",  x"21",  x"01",  x"fb",  x"cd",  x"1b",  x"55",  x"fd", -- 0198
         x"cb",  x"00",  x"46",  x"28",  x"0f",  x"21",  x"c0",  x"fb", -- 01A0
         x"cd",  x"1b",  x"55",  x"21",  x"81",  x"fc",  x"cd",  x"1b", -- 01A8
         x"55",  x"cd",  x"21",  x"59",  x"3a",  x"34",  x"0d",  x"3d", -- 01B0
         x"21",  x"3c",  x"0d",  x"b6",  x"ca",  x"f5",  x"53",  x"3a", -- 01B8
         x"49",  x"0d",  x"fe",  x"00",  x"28",  x"2d",  x"fa",  x"ea", -- 01C0
         x"51",  x"21",  x"4a",  x"0d",  x"35",  x"28",  x"21",  x"7e", -- 01C8
         x"e6",  x"07",  x"20",  x"1f",  x"3a",  x"49",  x"0d",  x"3d", -- 01D0
         x"32",  x"49",  x"0d",  x"28",  x"13",  x"c5",  x"47",  x"0e", -- 01D8
         x"0c",  x"21",  x"86",  x"f9",  x"cd",  x"41",  x"59",  x"c1", -- 01E0
         x"18",  x"09",  x"21",  x"4a",  x"0d",  x"35",  x"20",  x"03", -- 01E8
         x"cd",  x"0b",  x"59",  x"21",  x"02",  x"0d",  x"06",  x"10", -- 01F0
         x"7e",  x"e6",  x"f0",  x"fe",  x"a0",  x"20",  x"04",  x"7e", -- 01F8
         x"d6",  x"10",  x"77",  x"23",  x"10",  x"f2",  x"06",  x"10", -- 0200
         x"7e",  x"e6",  x"f0",  x"fe",  x"90",  x"20",  x"04",  x"7e", -- 0208
         x"c6",  x"10",  x"77",  x"23",  x"10",  x"f2",  x"cd",  x"ab", -- 0210
         x"58",  x"21",  x"2a",  x"0d",  x"cd",  x"ab",  x"58",  x"3a", -- 0218
         x"bf",  x"0c",  x"b7",  x"20",  x"40",  x"3e",  x"4d",  x"32", -- 0220
         x"bf",  x"0c",  x"3a",  x"56",  x"0c",  x"fd",  x"cb",  x"00", -- 0228
         x"46",  x"20",  x"09",  x"fe",  x"f0",  x"30",  x"05",  x"3e", -- 0230
         x"ff",  x"32",  x"56",  x"0c",  x"3d",  x"fe",  x"30",  x"38", -- 0238
         x"24",  x"32",  x"56",  x"0c",  x"6f",  x"e6",  x"03",  x"20", -- 0240
         x"0f",  x"ed",  x"5f",  x"e6",  x"03",  x"28",  x"09",  x"3a", -- 0248
         x"49",  x"0d",  x"b7",  x"20",  x"03",  x"cd",  x"cd",  x"58", -- 0250
         x"7d",  x"21",  x"46",  x"0d",  x"36",  x"00",  x"37",  x"cb", -- 0258
         x"16",  x"d6",  x"60",  x"30",  x"f9",  x"21",  x"3c",  x"fb", -- 0260
         x"cd",  x"96",  x"55",  x"11",  x"02",  x"0d",  x"cd",  x"30", -- 0268
         x"54",  x"fd",  x"cb",  x"00",  x"46",  x"ca",  x"5e",  x"53", -- 0270
         x"30",  x"06",  x"11",  x"22",  x"0d",  x"cd",  x"03",  x"55", -- 0278
         x"21",  x"c0",  x"fb",  x"cd",  x"96",  x"55",  x"11",  x"12", -- 0280
         x"0d",  x"cd",  x"84",  x"54",  x"30",  x"06",  x"11",  x"02", -- 0288
         x"0d",  x"cd",  x"ec",  x"54",  x"21",  x"bc",  x"fc",  x"cd", -- 0290
         x"96",  x"55",  x"11",  x"22",  x"0d",  x"cd",  x"30",  x"54", -- 0298
         x"30",  x"20",  x"11",  x"12",  x"0d",  x"cd",  x"ec",  x"54", -- 02A0
         x"3a",  x"32",  x"0d",  x"3d",  x"3d",  x"f2",  x"b2",  x"52", -- 02A8
         x"3e",  x"0f",  x"32",  x"32",  x"0d",  x"3a",  x"33",  x"0d", -- 02B0
         x"3c",  x"3c",  x"fe",  x"10",  x"20",  x"01",  x"af",  x"32", -- 02B8
         x"33",  x"0d",  x"fd",  x"cb",  x"00",  x"46",  x"28",  x"24", -- 02C0
         x"dd",  x"cb",  x"01",  x"76",  x"28",  x"1e",  x"21",  x"af", -- 02C8
         x"fc",  x"ed",  x"5f",  x"e6",  x"1f",  x"3c",  x"4f",  x"06", -- 02D0
         x"00",  x"3e",  x"a0",  x"ed",  x"b9",  x"20",  x"0d",  x"dd", -- 02D8
         x"21",  x"11",  x"5c",  x"3e",  x"03",  x"32",  x"4b",  x"0d", -- 02E0
         x"23",  x"22",  x"47",  x"0d",  x"cd",  x"c5",  x"57",  x"3a", -- 02E8
         x"00",  x"0d",  x"3d",  x"20",  x"02",  x"3e",  x"02",  x"32", -- 02F0
         x"00",  x"0d",  x"cd",  x"96",  x"55",  x"fd",  x"cb",  x"00", -- 02F8
         x"46",  x"28",  x"67",  x"db",  x"84",  x"1f",  x"38",  x"4f", -- 0300
         x"3a",  x"3e",  x"0d",  x"b7",  x"c2",  x"b4",  x"51",  x"3c", -- 0308
         x"32",  x"3e",  x"0d",  x"3a",  x"34",  x"0d",  x"fe",  x"01", -- 0310
         x"c2",  x"b4",  x"51",  x"21",  x"3c",  x"0d",  x"35",  x"fa", -- 0318
         x"f5",  x"53",  x"cd",  x"21",  x"59",  x"3e",  x"1c",  x"32", -- 0320
         x"34",  x"0d",  x"3a",  x"35",  x"0d",  x"32",  x"36",  x"0d", -- 0328
         x"3e",  x"20",  x"32",  x"3b",  x"0d",  x"2a",  x"39",  x"0d", -- 0330
         x"01",  x"c1",  x"ff",  x"09",  x"3a",  x"35",  x"0d",  x"77", -- 0338
         x"22",  x"37",  x"0d",  x"21",  x"47",  x"5c",  x"7e",  x"32", -- 0340
         x"60",  x"0c",  x"23",  x"7e",  x"32",  x"61",  x"0c",  x"3e", -- 0348
         x"55",  x"32",  x"5a",  x"0c",  x"c3",  x"b4",  x"51",  x"af", -- 0350
         x"32",  x"3e",  x"0d",  x"c3",  x"b4",  x"51",  x"d2",  x"c2", -- 0358
         x"52",  x"11",  x"02",  x"0d",  x"cd",  x"03",  x"55",  x"c3", -- 0360
         x"a8",  x"52",  x"11",  x"92",  x"ff",  x"21",  x"0a",  x"03", -- 0368
         x"01",  x"1b",  x"00",  x"ed",  x"b0",  x"cd",  x"c7",  x"01", -- 0370
         x"cd",  x"c7",  x"01",  x"cd",  x"6f",  x"57",  x"21",  x"83", -- 0378
         x"fc",  x"3e",  x"a0",  x"cd",  x"79",  x"55",  x"21",  x"43", -- 0380
         x"fd",  x"3e",  x"80",  x"cd",  x"79",  x"55",  x"21",  x"03", -- 0388
         x"fe",  x"3e",  x"b0",  x"cd",  x"79",  x"55",  x"06",  x"08", -- 0390
         x"21",  x"9b",  x"5a",  x"c5",  x"cd",  x"13",  x"57",  x"c1", -- 0398
         x"10",  x"f9",  x"21",  x"a1",  x"fc",  x"36",  x"d0",  x"23", -- 03A0
         x"36",  x"d0",  x"21",  x"21",  x"fd",  x"36",  x"d8",  x"23", -- 03A8
         x"36",  x"d8",  x"23",  x"23",  x"23",  x"36",  x"2d",  x"21", -- 03B0
         x"a1",  x"fd",  x"36",  x"d6",  x"23",  x"36",  x"d6",  x"23", -- 03B8
         x"23",  x"23",  x"36",  x"2d",  x"21",  x"21",  x"fe",  x"36", -- 03C0
         x"da",  x"23",  x"36",  x"da",  x"23",  x"23",  x"23",  x"36", -- 03C8
         x"2d",  x"cd",  x"9a",  x"01",  x"c2",  x"f1",  x"00",  x"3a", -- 03D0
         x"03",  x"0c",  x"b7",  x"ca",  x"b4",  x"51",  x"fd",  x"36", -- 03D8
         x"00",  x"ff",  x"cd",  x"26",  x"03",  x"2a",  x"00",  x"0c", -- 03E0
         x"23",  x"22",  x"00",  x"0c",  x"21",  x"00",  x"00",  x"22", -- 03E8
         x"18",  x"0c",  x"c3",  x"45",  x"50",  x"af",  x"32",  x"03", -- 03F0
         x"0c",  x"fd",  x"77",  x"00",  x"21",  x"00",  x"fb",  x"36"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
