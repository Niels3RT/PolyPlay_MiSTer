library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom2_1400 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom2_1400;

architecture rtl of rom2_1400 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"49",  x"4e",  x"45",  x"4e",  x"20",  x"50",  x"52",  x"4f", -- 0000
         x"42",  x"45",  x"4c",  x"41",  x"55",  x"46",  x"20",  x"20", -- 0008
         x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20", -- 0010
         x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20", -- 0018
         x"90",  x"fc",  x"1d",  x"4d",  x"49",  x"54",  x"20",  x"56", -- 0020
         x"45",  x"52",  x"47",  x"52",  x"4f",  x"45",  x"53",  x"53", -- 0028
         x"45",  x"52",  x"54",  x"45",  x"52",  x"20",  x"54",  x"4f", -- 0030
         x"52",  x"57",  x"45",  x"49",  x"54",  x"45",  x"20",  x"3f", -- 0038
         x"98",  x"fd",  x"1e",  x"4a",  x"41",  x"20",  x"3c",  x"2d", -- 0040
         x"2d",  x"20",  x"53",  x"54",  x"45",  x"55",  x"45",  x"52", -- 0048
         x"4b",  x"4e",  x"55",  x"45",  x"50",  x"50",  x"45",  x"4c", -- 0050
         x"20",  x"2d",  x"2d",  x"3e",  x"20",  x"4e",  x"45",  x"49", -- 0058
         x"4e",  x"50",  x"f9",  x"19",  x"2a",  x"2a",  x"20",  x"44", -- 0060
         x"49",  x"53",  x"51",  x"55",  x"41",  x"4c",  x"49",  x"46", -- 0068
         x"49",  x"4b",  x"41",  x"54",  x"49",  x"4f",  x"4e",  x"20", -- 0070
         x"4e",  x"41",  x"43",  x"48",  x"3a",  x"6d",  x"f9",  x"0a", -- 0078
         x"20",  x"4d",  x"45",  x"54",  x"45",  x"52",  x"4e",  x"20", -- 0080
         x"2a",  x"2a",  x"84",  x"f8",  x"05",  x"2e",  x"4c",  x"41", -- 0088
         x"55",  x"46",  x"04",  x"fb",  x"06",  x"20",  x"4c",  x"41", -- 0090
         x"55",  x"46",  x"20",  x"0b",  x"fb",  x"0e",  x"20",  x"20", -- 0098
         x"20",  x"54",  x"4f",  x"52",  x"57",  x"45",  x"49",  x"54", -- 00A0
         x"45",  x"20",  x"20",  x"20",  x"1a",  x"fb",  x"12",  x"20", -- 00A8
         x"20",  x"20",  x"20",  x"20",  x"46",  x"41",  x"48",  x"52", -- 00B0
         x"5a",  x"45",  x"49",  x"54",  x"20",  x"20",  x"20",  x"20", -- 00B8
         x"20",  x"2d",  x"fb",  x"0f",  x"20",  x"20",  x"20",  x"42", -- 00C0
         x"45",  x"57",  x"45",  x"52",  x"54",  x"55",  x"4e",  x"47", -- 00C8
         x"20",  x"20",  x"20",  x"d4",  x"ff",  x"18",  x"2a",  x"2a", -- 00D0
         x"2a",  x"20",  x"45",  x"4e",  x"44",  x"45",  x"20",  x"44", -- 00D8
         x"45",  x"53",  x"20",  x"53",  x"50",  x"49",  x"45",  x"4c", -- 00E0
         x"45",  x"53",  x"20",  x"2a",  x"2a",  x"2a",  x"d0",  x"fe", -- 00E8
         x"20",  x"53",  x"20",  x"49",  x"20",  x"4e",  x"20",  x"44", -- 00F0
         x"20",  x"20",  x"20",  x"53",  x"20",  x"49",  x"20",  x"45", -- 00F8
         x"20",  x"20",  x"20",  x"42",  x"20",  x"45",  x"20",  x"53", -- 0100
         x"20",  x"53",  x"20",  x"45",  x"20",  x"52",  x"20",  x"20", -- 0108
         x"3f",  x"ac",  x"f8",  x"09",  x"54",  x"4f",  x"52",  x"57", -- 0110
         x"45",  x"49",  x"54",  x"45",  x"3a",  x"06",  x"20",  x"4d", -- 0118
         x"45",  x"54",  x"45",  x"52",  x"09",  x"20",  x"53",  x"45", -- 0120
         x"4b",  x"55",  x"4e",  x"44",  x"45",  x"4e",  x"07",  x"20", -- 0128
         x"50",  x"55",  x"4e",  x"4b",  x"54",  x"45",  x"0d",  x"41", -- 0130
         x"55",  x"53",  x"47",  x"45",  x"53",  x"43",  x"48",  x"49", -- 0138
         x"45",  x"44",  x"45",  x"4e",  x"08",  x"80",  x"02",  x"60", -- 0140
         x"00",  x"3f",  x"ff",  x"02",  x"40",  x"44",  x"80",  x"00", -- 0148
         x"3f",  x"ff",  x"00",  x"10",  x"00",  x"82",  x"01",  x"18", -- 0150
         x"9c",  x"82",  x"01",  x"08",  x"d0",  x"82",  x"01",  x"10", -- 0158
         x"af",  x"82",  x"01",  x"10",  x"c4",  x"82",  x"01",  x"20", -- 0160
         x"00",  x"98",  x"01",  x"10",  x"00",  x"82",  x"01",  x"18", -- 0168
         x"00",  x"82",  x"01",  x"48",  x"14",  x"82",  x"01",  x"10", -- 0170
         x"e9",  x"82",  x"01",  x"50",  x"14",  x"82",  x"01",  x"60", -- 0178
         x"12",  x"00",  x"20",  x"c4",  x"82",  x"01",  x"20",  x"93", -- 0180
         x"82",  x"01",  x"58",  x"12",  x"82",  x"01",  x"48",  x"12", -- 0188
         x"82",  x"01",  x"58",  x"12",  x"98",  x"01",  x"10",  x"c4", -- 0190
         x"82",  x"01",  x"18",  x"e9",  x"82",  x"01",  x"10",  x"c4", -- 0198
         x"82",  x"01",  x"3f",  x"93",  x"18",  x"93",  x"82",  x"01", -- 01A0
         x"08",  x"9c",  x"82",  x"01",  x"18",  x"af",  x"82",  x"01", -- 01A8
         x"08",  x"e9",  x"82",  x"01",  x"3f",  x"c4",  x"82",  x"01", -- 01B0
         x"18",  x"dc",  x"82",  x"01",  x"08",  x"dc",  x"82",  x"01", -- 01B8
         x"18",  x"c4",  x"82",  x"01",  x"08",  x"af",  x"82",  x"01", -- 01C0
         x"3f",  x"9c",  x"18",  x"9c",  x"82",  x"01",  x"08",  x"af", -- 01C8
         x"82",  x"01",  x"18",  x"c4",  x"82",  x"01",  x"08",  x"dc", -- 01D0
         x"82",  x"01",  x"3f",  x"e9",  x"18",  x"e9",  x"8f",  x"01", -- 01D8
         x"00",  x"8f",  x"01",  x"48",  x"12",  x"82",  x"01",  x"08", -- 01E0
         x"e9",  x"82",  x"01",  x"08",  x"c4",  x"82",  x"01",  x"20", -- 01E8
         x"93",  x"00",  x"08",  x"00",  x"0d",  x"18",  x"3c",  x"7e", -- 01F0
         x"ff",  x"ff",  x"7e",  x"3c",  x"18",  x"00",  x"00",  x"00", -- 01F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"36",  x"0d",  x"03", -- 0200
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"80",  x"60", -- 0208
         x"d8",  x"36",  x"0d",  x"03",  x"00",  x"00",  x"00",  x"00", -- 0210
         x"00",  x"00",  x"80",  x"60",  x"d8",  x"0d",  x"06",  x"01", -- 0218
         x"00",  x"00",  x"00",  x"00",  x"00",  x"80",  x"c0",  x"b0", -- 0220
         x"d8",  x"36",  x"1b",  x"06",  x"03",  x"00",  x"00",  x"00", -- 0228
         x"00",  x"00",  x"00",  x"c0",  x"60",  x"03",  x"01",  x"00", -- 0230
         x"00",  x"00",  x"00",  x"00",  x"00",  x"60",  x"b0",  x"d8", -- 0238
         x"6c",  x"36",  x"1b",  x"0d",  x"06",  x"00",  x"00",  x"00", -- 0240
         x"00",  x"00",  x"00",  x"80",  x"c0",  x"00",  x"00",  x"00", -- 0248
         x"00",  x"00",  x"00",  x"00",  x"00",  x"90",  x"d8",  x"48", -- 0250
         x"6c",  x"24",  x"36",  x"12",  x"1b",  x"10",  x"00",  x"01", -- 0258
         x"24",  x"24",  x"24",  x"24",  x"24",  x"24",  x"24",  x"24", -- 0260
         x"08",  x"00",  x"0c",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0268
         x"00",  x"00",  x"00",  x"09",  x"1b",  x"12",  x"36",  x"24", -- 0270
         x"6c",  x"48",  x"d8",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0278
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0280
         x"00",  x"01",  x"03",  x"06",  x"0d",  x"1b",  x"36",  x"6c", -- 0288
         x"d8",  x"b0",  x"60",  x"c0",  x"80",  x"00",  x"00",  x"00", -- 0290
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0298
         x"00",  x"03",  x"06",  x"01",  x"03",  x"0d",  x"1b",  x"6c", -- 02A0
         x"d8",  x"60",  x"c0",  x"b0",  x"60",  x"80",  x"00",  x"00", -- 02A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02B0
         x"01",  x"06",  x"1b",  x"00",  x"01",  x"06",  x"1b",  x"6c", -- 02B8
         x"b0",  x"c0",  x"00",  x"6c",  x"b0",  x"c0",  x"00",  x"00", -- 02C0
         x"00",  x"00",  x"00",  x"08",  x"00",  x"07",  x"ff",  x"ff", -- 02C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"00", -- 02D0
         x"00",  x"00",  x"00",  x"00",  x"03",  x"07",  x"3c",  x"7e", -- 02D8
         x"7e",  x"00",  x"00",  x"3c",  x"ff",  x"ff",  x"00",  x"00", -- 02E0
         x"00",  x"00",  x"00",  x"00",  x"c0",  x"e0",  x"07",  x"cd", -- 02E8
         x"79",  x"31",  x"01",  x"01",  x"01",  x"01",  x"ff",  x"cb", -- 02F0
         x"c3",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"e0",  x"b3", -- 02F8
         x"be",  x"9c",  x"80",  x"80",  x"80",  x"80",  x"18",  x"00", -- 0300
         x"02",  x"01",  x"03",  x"07",  x"0f",  x"1e",  x"1e",  x"0e", -- 0308
         x"07",  x"ff",  x"fe",  x"bc",  x"78",  x"78",  x"f0",  x"70", -- 0310
         x"38",  x"10",  x"00",  x"02",  x"03",  x"01",  x"00",  x"00", -- 0318
         x"00",  x"00",  x"00",  x"00",  x"38",  x"9c",  x"da",  x"00", -- 0320
         x"00",  x"00",  x"00",  x"00",  x"20",  x"00",  x"02",  x"01", -- 0328
         x"03",  x"07",  x"0f",  x"1e",  x"1e",  x"07",  x"03",  x"ff", -- 0330
         x"fe",  x"bc",  x"78",  x"78",  x"f0",  x"38",  x"1c",  x"10", -- 0338
         x"00",  x"02",  x"01",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0340
         x"00",  x"00",  x"1c",  x"c6",  x"66",  x"00",  x"00",  x"00", -- 0348
         x"00",  x"00",  x"20",  x"00",  x"03",  x"01",  x"01",  x"00", -- 0350
         x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"f7", -- 0358
         x"e7",  x"f7",  x"e7",  x"e7",  x"66",  x"80",  x"80",  x"00", -- 0360
         x"00",  x"00",  x"00",  x"00",  x"00",  x"10",  x"00",  x"01", -- 0368
         x"66",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"24", -- 0370
         x"28",  x"00",  x"02",  x"ff",  x"7f",  x"3d",  x"1e",  x"1e", -- 0378
         x"0f",  x"1c",  x"39",  x"80",  x"c0",  x"e0",  x"f0",  x"78", -- 0380
         x"78",  x"e0",  x"c0",  x"10",  x"00",  x"02",  x"39",  x"73", -- 0388
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"80",  x"00", -- 0390
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"20",  x"00", -- 0398
         x"02",  x"ff",  x"7f",  x"3d",  x"1e",  x"1e",  x"0f",  x"0e", -- 03A0
         x"1c",  x"80",  x"c0",  x"e0",  x"f0",  x"78",  x"78",  x"70", -- 03A8
         x"e0",  x"10",  x"00",  x"05",  x"70",  x"39",  x"e3",  x"00", -- 03B0
         x"00",  x"00",  x"00",  x"00",  x"c0",  x"80",  x"00",  x"00", -- 03B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03C0
         x"00",  x"00",  x"00",  x"00",  x"07",  x"0f",  x"80",  x"81", -- 03C8
         x"86",  x"9e",  x"b0",  x"b0",  x"e0",  x"f0",  x"01",  x"e1", -- 03D0
         x"39",  x"3d",  x"07",  x"07",  x"10",  x"00",  x"02",  x"30", -- 03D8
         x"1e",  x"0e",  x"07",  x"00",  x"00",  x"00",  x"00",  x"06", -- 03E0
         x"3c",  x"3c",  x"f0",  x"00",  x"00",  x"00",  x"00",  x"08", -- 03E8
         x"01",  x"03",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff", -- 03F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"18",  x"18",  x"00"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
