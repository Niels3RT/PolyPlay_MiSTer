library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_6000 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_6000;

architecture rtl of rom1_6000 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"cd",  x"b7",  x"01",  x"cd",  x"b7",  x"02",  x"11",  x"00", -- 0000
         x"ec",  x"21",  x"21",  x"6a",  x"3a",  x"f3",  x"72",  x"47", -- 0008
         x"c5",  x"4e",  x"23",  x"46",  x"23",  x"7e",  x"23",  x"eb", -- 0010
         x"09",  x"eb",  x"47",  x"c5",  x"01",  x"08",  x"00",  x"ed", -- 0018
         x"b0",  x"c1",  x"10",  x"f7",  x"c1",  x"10",  x"e9",  x"fd", -- 0020
         x"21",  x"2e",  x"0d",  x"fd",  x"36",  x"00",  x"00",  x"3e", -- 0028
         x"03",  x"32",  x"2d",  x"0d",  x"21",  x"00",  x"f8",  x"11", -- 0030
         x"01",  x"f8",  x"01",  x"ff",  x"07",  x"36",  x"20",  x"ed", -- 0038
         x"b0",  x"dd",  x"21",  x"01",  x"0d",  x"dd",  x"36",  x"00", -- 0040
         x"80",  x"dd",  x"36",  x"01",  x"00",  x"dd",  x"36",  x"02", -- 0048
         x"04",  x"dd",  x"36",  x"03",  x"10",  x"dd",  x"36",  x"04", -- 0050
         x"10",  x"dd",  x"36",  x"07",  x"07",  x"dd",  x"21",  x"09", -- 0058
         x"0d",  x"dd",  x"36",  x"00",  x"80",  x"dd",  x"36",  x"01", -- 0060
         x"00",  x"dd",  x"36",  x"02",  x"04",  x"dd",  x"36",  x"03", -- 0068
         x"28",  x"dd",  x"36",  x"04",  x"28",  x"dd",  x"36",  x"07", -- 0070
         x"07",  x"dd",  x"36",  x"08",  x"00",  x"af",  x"32",  x"00", -- 0078
         x"0d",  x"32",  x"2b",  x"0d",  x"32",  x"2c",  x"0d",  x"32", -- 0080
         x"56",  x"0c",  x"32",  x"33",  x"0d",  x"21",  x"00",  x"00", -- 0088
         x"22",  x"13",  x"0d",  x"22",  x"2f",  x"0d",  x"3e",  x"fd", -- 0090
         x"32",  x"15",  x"0d",  x"cd",  x"49",  x"66",  x"06",  x"40", -- 0098
         x"21",  x"40",  x"f8",  x"3e",  x"fc",  x"77",  x"23",  x"10", -- 00A0
         x"fc",  x"cd",  x"72",  x"66",  x"2e",  x"67",  x"21",  x"0c", -- 00A8
         x"f8",  x"22",  x"3f",  x"0c",  x"2a",  x"10",  x"0c",  x"22", -- 00B0
         x"3d",  x"0c",  x"cd",  x"70",  x"02",  x"21",  x"1e",  x"f8", -- 00B8
         x"22",  x"3f",  x"0c",  x"2a",  x"18",  x"0c",  x"22",  x"3d", -- 00C0
         x"0c",  x"cd",  x"70",  x"02",  x"fd",  x"cb",  x"00",  x"46", -- 00C8
         x"20",  x"69",  x"11",  x"92",  x"ff",  x"21",  x"0a",  x"03", -- 00D0
         x"01",  x"1b",  x"00",  x"ed",  x"b0",  x"06",  x"05",  x"21", -- 00D8
         x"cc",  x"67",  x"c5",  x"cd",  x"7a",  x"66",  x"c1",  x"10", -- 00E0
         x"f9",  x"06",  x"1d",  x"3e",  x"ff",  x"21",  x"90",  x"f9", -- 00E8
         x"77",  x"23",  x"10",  x"fc",  x"06",  x"40",  x"3e",  x"80", -- 00F0
         x"21",  x"40",  x"fe",  x"77",  x"23",  x"10",  x"fc",  x"21", -- 00F8
         x"43",  x"fa",  x"dd",  x"21",  x"01",  x"0d",  x"af",  x"32", -- 0100
         x"16",  x"0d",  x"cd",  x"7f",  x"65",  x"21",  x"83",  x"fb", -- 0108
         x"dd",  x"21",  x"09",  x"0d",  x"3e",  x"01",  x"32",  x"16", -- 0110
         x"0d",  x"cd",  x"7f",  x"65",  x"cd",  x"9a",  x"01",  x"c2", -- 0118
         x"f1",  x"00",  x"3a",  x"03",  x"0c",  x"b7",  x"28",  x"f4", -- 0120
         x"21",  x"f4",  x"69",  x"cd",  x"e0",  x"01",  x"21",  x"00", -- 0128
         x"00",  x"22",  x"18",  x"0c",  x"fd",  x"36",  x"00",  x"01", -- 0130
         x"c3",  x"34",  x"60",  x"cd",  x"72",  x"66",  x"b7",  x"67", -- 0138
         x"21",  x"2d",  x"0d",  x"cb",  x"4e",  x"20",  x"05",  x"21", -- 0140
         x"d2",  x"f8",  x"36",  x"32",  x"cd",  x"72",  x"66",  x"c2", -- 0148
         x"67",  x"dd",  x"21",  x"74",  x"69",  x"0e",  x"fd",  x"21", -- 0150
         x"c9",  x"f8",  x"cd",  x"90",  x"66",  x"21",  x"f7",  x"f8", -- 0158
         x"cd",  x"90",  x"66",  x"21",  x"a5",  x"fa",  x"cd",  x"90", -- 0160
         x"66",  x"21",  x"77",  x"fc",  x"cd",  x"90",  x"66",  x"21", -- 0168
         x"e1",  x"ff",  x"cd",  x"90",  x"66",  x"21",  x"2d",  x"0d", -- 0170
         x"cb",  x"46",  x"20",  x"06",  x"21",  x"ce",  x"f9",  x"cd", -- 0178
         x"90",  x"66",  x"dd",  x"21",  x"23",  x"69",  x"21",  x"c1", -- 0180
         x"f8",  x"0e",  x"ff",  x"cd",  x"90",  x"66",  x"21",  x"b7", -- 0188
         x"fa",  x"cd",  x"90",  x"66",  x"21",  x"ca",  x"fa",  x"cd", -- 0190
         x"90",  x"66",  x"dd",  x"21",  x"5c",  x"69",  x"0e",  x"fe", -- 0198
         x"21",  x"50",  x"fc",  x"cd",  x"90",  x"66",  x"dd",  x"21", -- 01A0
         x"6e",  x"69",  x"21",  x"5a",  x"fc",  x"cd",  x"90",  x"66", -- 01A8
         x"0e",  x"fa",  x"cd",  x"d4",  x"66",  x"21",  x"2d",  x"0d", -- 01B0
         x"cb",  x"46",  x"20",  x"17",  x"21",  x"46",  x"fc",  x"22", -- 01B8
         x"0e",  x"0d",  x"dd",  x"21",  x"09",  x"0d",  x"3e",  x"01", -- 01C0
         x"32",  x"16",  x"0d",  x"cd",  x"7f",  x"65",  x"21",  x"41", -- 01C8
         x"fc",  x"18",  x"15",  x"21",  x"41",  x"fc",  x"22",  x"0e", -- 01D0
         x"0d",  x"dd",  x"21",  x"09",  x"0d",  x"3e",  x"01",  x"32", -- 01D8
         x"16",  x"0d",  x"cd",  x"7f",  x"65",  x"21",  x"45",  x"fc", -- 01E0
         x"22",  x"06",  x"0d",  x"dd",  x"21",  x"01",  x"0d",  x"af", -- 01E8
         x"32",  x"16",  x"0d",  x"cd",  x"7f",  x"65",  x"e5",  x"21", -- 01F0
         x"fc",  x"68",  x"cd",  x"e0",  x"01",  x"e1",  x"3e",  x"4d", -- 01F8
         x"32",  x"bf",  x"0c",  x"e5",  x"af",  x"32",  x"00",  x"0d", -- 0200
         x"3a",  x"16",  x"0d",  x"b7",  x"20",  x"0f",  x"3e",  x"09", -- 0208
         x"dd",  x"96",  x"07",  x"cb",  x"3f",  x"f6",  x"30",  x"21", -- 0210
         x"52",  x"f9",  x"77",  x"e1",  x"e5",  x"dd",  x"e5",  x"7c", -- 0218
         x"e6",  x"07",  x"fe",  x"04",  x"c2",  x"bc",  x"62",  x"7d", -- 0220
         x"fe",  x"09",  x"30",  x"43",  x"dd",  x"cb",  x"07",  x"46", -- 0228
         x"c2",  x"bc",  x"62",  x"dd",  x"35",  x"07",  x"fa",  x"6c", -- 0230
         x"64",  x"21",  x"2b",  x"0d",  x"35",  x"cb",  x"46",  x"20", -- 0238
         x"7b",  x"cd",  x"06",  x"67",  x"21",  x"50",  x"fc",  x"e5", -- 0240
         x"0e",  x"fe",  x"dd",  x"7e",  x"02",  x"fe",  x"08",  x"30", -- 0248
         x"0f",  x"dd",  x"21",  x"5c",  x"69",  x"cd",  x"90",  x"66", -- 0250
         x"e1",  x"0e",  x"20",  x"cd",  x"90",  x"66",  x"18",  x"5c", -- 0258
         x"dd",  x"21",  x"62",  x"69",  x"cd",  x"90",  x"66",  x"e1", -- 0260
         x"0e",  x"20",  x"cd",  x"90",  x"66",  x"18",  x"4d",  x"d6", -- 0268
         x"5b",  x"fe",  x"08",  x"30",  x"47",  x"dd",  x"cb",  x"07", -- 0270
         x"46",  x"28",  x"41",  x"dd",  x"35",  x"07",  x"0e",  x"20", -- 0278
         x"20",  x"02",  x"0e",  x"fb",  x"cd",  x"d4",  x"66",  x"21", -- 0280
         x"2c",  x"0d",  x"35",  x"cb",  x"46",  x"20",  x"2d",  x"cd", -- 0288
         x"06",  x"67",  x"21",  x"5a",  x"fc",  x"e5",  x"0e",  x"fe", -- 0290
         x"dd",  x"7e",  x"02",  x"3d",  x"fe",  x"08",  x"30",  x"0f", -- 0298
         x"dd",  x"21",  x"68",  x"69",  x"cd",  x"90",  x"66",  x"e1", -- 02A0
         x"0e",  x"20",  x"cd",  x"90",  x"66",  x"18",  x"0d",  x"dd", -- 02A8
         x"21",  x"6e",  x"69",  x"cd",  x"90",  x"66",  x"e1",  x"0e", -- 02B0
         x"20",  x"cd",  x"90",  x"66",  x"dd",  x"e1",  x"dd",  x"7e", -- 02B8
         x"03",  x"21",  x"12",  x"0d",  x"34",  x"cb",  x"46",  x"20", -- 02C0
         x"0f",  x"c6",  x"bd",  x"32",  x"60",  x"0c",  x"3c",  x"3c", -- 02C8
         x"32",  x"61",  x"0c",  x"3e",  x"55",  x"32",  x"5a",  x"0c", -- 02D0
         x"e1",  x"dd",  x"75",  x"05",  x"dd",  x"74",  x"06",  x"3e", -- 02D8
         x"b0",  x"3d",  x"20",  x"fd",  x"3a",  x"bf",  x"0c",  x"b7", -- 02E0
         x"20",  x"27",  x"3e",  x"4d",  x"32",  x"bf",  x"0c",  x"3a", -- 02E8
         x"13",  x"0d",  x"3c",  x"fe",  x"64",  x"d2",  x"4a",  x"65", -- 02F0
         x"32",  x"13",  x"0d",  x"32",  x"3d",  x"0c",  x"e5",  x"21", -- 02F8
         x"2d",  x"f8",  x"22",  x"3f",  x"0c",  x"cd",  x"70",  x"02", -- 0300
         x"36",  x"20",  x"2b",  x"36",  x"20",  x"2b",  x"36",  x"2c", -- 0308
         x"e1",  x"dd",  x"21",  x"01",  x"0d",  x"dd",  x"35",  x"04", -- 0310
         x"28",  x"4c",  x"dd",  x"21",  x"09",  x"0d",  x"dd",  x"35", -- 0318
         x"04",  x"20",  x"bc",  x"3a",  x"08",  x"0d",  x"dd",  x"96", -- 0320
         x"07",  x"30",  x"0c",  x"dd",  x"35",  x"03",  x"dd",  x"35", -- 0328
         x"03",  x"dd",  x"36",  x"08",  x"fc",  x"18",  x"06",  x"28", -- 0330
         x"04",  x"dd",  x"36",  x"08",  x"02",  x"3a",  x"04",  x"0d", -- 0338
         x"dd",  x"86",  x"03",  x"dd",  x"86",  x"03",  x"dd",  x"86", -- 0340
         x"03",  x"cb",  x"3f",  x"cb",  x"3f",  x"dd",  x"77",  x"03", -- 0348
         x"dd",  x"86",  x"08",  x"dd",  x"77",  x"04",  x"3e",  x"01", -- 0350
         x"32",  x"16",  x"0d",  x"2a",  x"0e",  x"0d",  x"3e",  x"fc", -- 0358
         x"32",  x"15",  x"0d",  x"e5",  x"18",  x"4a",  x"dd",  x"7e", -- 0360
         x"03",  x"dd",  x"77",  x"04",  x"af",  x"32",  x"16",  x"0d", -- 0368
         x"2a",  x"06",  x"0d",  x"3e",  x"fd",  x"32",  x"15",  x"0d", -- 0370
         x"db",  x"84",  x"cb",  x"47",  x"4f",  x"20",  x"10",  x"3e", -- 0378
         x"10",  x"06",  x"04",  x"dd",  x"35",  x"03",  x"dd",  x"be", -- 0380
         x"03",  x"30",  x"04",  x"10",  x"f6",  x"18",  x"0d",  x"3e", -- 0388
         x"40",  x"dd",  x"34",  x"03",  x"dd",  x"be",  x"03",  x"30", -- 0390
         x"03",  x"dd",  x"35",  x"03",  x"79",  x"e5",  x"e6",  x"1e", -- 0398
         x"21",  x"ec",  x"69",  x"01",  x"08",  x"00",  x"ed",  x"b1", -- 03A0
         x"c2",  x"53",  x"64",  x"cb",  x"21",  x"dd",  x"71",  x"02", -- 03A8
         x"3e",  x"38",  x"dd",  x"ae",  x"01",  x"dd",  x"77",  x"01", -- 03B0
         x"cd",  x"e3",  x"66",  x"c2",  x"53",  x"64",  x"dd",  x"7e", -- 03B8
         x"02",  x"cd",  x"c8",  x"66",  x"e1",  x"cd",  x"f8",  x"65", -- 03C0
         x"cd",  x"01",  x"66",  x"19",  x"cd",  x"3f",  x"66",  x"3a", -- 03C8
         x"00",  x"0d",  x"b7",  x"28",  x"7f",  x"cb",  x"7f",  x"c2", -- 03D0
         x"64",  x"64",  x"ed",  x"52",  x"e5",  x"06",  x"05",  x"cd", -- 03D8
         x"63",  x"66",  x"10",  x"fb",  x"21",  x"00",  x"0d",  x"36", -- 03E0
         x"00",  x"dd",  x"7e",  x"02",  x"3d",  x"3d",  x"e6",  x"0e", -- 03E8
         x"dd",  x"77",  x"02",  x"cd",  x"c8",  x"66",  x"cd",  x"de", -- 03F0
         x"66",  x"e1",  x"19",  x"cd",  x"3f",  x"66",  x"3a",  x"00"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
