library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom2_1000 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom2_1000;

architecture rtl of rom2_1000 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"cd",  x"b7",  x"01",  x"cd",  x"b7",  x"02",  x"fd",  x"21", -- 0000
         x"56",  x"0d",  x"11",  x"00",  x"ec",  x"21",  x"f2",  x"15", -- 0008
         x"3a",  x"ad",  x"1b",  x"47",  x"c5",  x"4e",  x"23",  x"46", -- 0010
         x"23",  x"7e",  x"23",  x"eb",  x"09",  x"eb",  x"47",  x"c5", -- 0018
         x"01",  x"08",  x"00",  x"ed",  x"b0",  x"c1",  x"10",  x"f7", -- 0020
         x"c1",  x"10",  x"e9",  x"11",  x"18",  x"f0",  x"21",  x"05", -- 0028
         x"16",  x"01",  x"58",  x"00",  x"ed",  x"b0",  x"23",  x"23", -- 0030
         x"23",  x"11",  x"80",  x"f0",  x"01",  x"08",  x"00",  x"ed", -- 0038
         x"b0",  x"23",  x"23",  x"23",  x"11",  x"90",  x"f0",  x"01", -- 0040
         x"60",  x"00",  x"ed",  x"b0",  x"cd",  x"9a",  x"01",  x"c2", -- 0048
         x"f1",  x"00",  x"3a",  x"03",  x"0c",  x"b7",  x"20",  x"1b", -- 0050
         x"11",  x"92",  x"ff",  x"21",  x"0a",  x"03",  x"01",  x"1b", -- 0058
         x"00",  x"ed",  x"b0",  x"cd",  x"f0",  x"05",  x"ee",  x"14", -- 0060
         x"21",  x"00",  x"fe",  x"3e",  x"80",  x"06",  x"40",  x"77", -- 0068
         x"23",  x"10",  x"fc",  x"af",  x"21",  x"57",  x"0d",  x"01", -- 0070
         x"00",  x"0d",  x"c5",  x"ed",  x"42",  x"e5",  x"c1",  x"e1", -- 0078
         x"11",  x"01",  x"0d",  x"77",  x"ed",  x"b0",  x"3a",  x"03", -- 0080
         x"0c",  x"fd",  x"77",  x"00",  x"21",  x"1a",  x"0d",  x"36", -- 0088
         x"0f",  x"dd",  x"21",  x"1d",  x"0d",  x"cd",  x"f0",  x"05", -- 0090
         x"ae",  x"13",  x"21",  x"0b",  x"f8",  x"22",  x"3f",  x"0c", -- 0098
         x"2a",  x"0e",  x"0c",  x"22",  x"3d",  x"0c",  x"cd",  x"70", -- 00A0
         x"02",  x"21",  x"40",  x"f8",  x"06",  x"40",  x"36",  x"9f", -- 00A8
         x"23",  x"10",  x"fb",  x"fd",  x"cb",  x"00",  x"46",  x"28", -- 00B0
         x"36",  x"21",  x"01",  x"80",  x"22",  x"57",  x"0d",  x"21", -- 00B8
         x"53",  x"15",  x"cd",  x"d4",  x"01",  x"2a",  x"00",  x"0c", -- 00C0
         x"23",  x"22",  x"00",  x"0c",  x"3e",  x"1e",  x"21",  x"80", -- 00C8
         x"f8",  x"cd",  x"bc",  x"01",  x"06",  x"03",  x"21",  x"ee", -- 00D0
         x"13",  x"c5",  x"cd",  x"f8",  x"05",  x"c1",  x"10",  x"f9", -- 00D8
         x"db",  x"84",  x"cb",  x"4f",  x"28",  x"09",  x"cb",  x"57", -- 00E0
         x"20",  x"f6",  x"21",  x"1a",  x"0d",  x"cb",  x"26",  x"21", -- 00E8
         x"07",  x"0d",  x"34",  x"3e",  x"06",  x"be",  x"d2",  x"0e", -- 00F0
         x"11",  x"af",  x"32",  x"03",  x"0c",  x"fd",  x"77",  x"00", -- 00F8
         x"cd",  x"f0",  x"05",  x"d3",  x"14",  x"21",  x"82",  x"15", -- 0100
         x"cd",  x"e0",  x"01",  x"c3",  x"f1",  x"00",  x"21",  x"d8", -- 0108
         x"ff",  x"fd",  x"cb",  x"00",  x"46",  x"20",  x"02",  x"25", -- 0110
         x"25",  x"22",  x"01",  x"0d",  x"21",  x"08",  x"0d",  x"36", -- 0118
         x"82",  x"21",  x"09",  x"0d",  x"36",  x"01",  x"af",  x"32", -- 0120
         x"05",  x"0d",  x"32",  x"00",  x"0d",  x"32",  x"06",  x"0d", -- 0128
         x"3e",  x"07",  x"32",  x"04",  x"0d",  x"3e",  x"4d",  x"32", -- 0130
         x"bf",  x"0c",  x"3e",  x"90",  x"32",  x"56",  x"0c",  x"cd", -- 0138
         x"d8",  x"06",  x"21",  x"82",  x"f8",  x"22",  x"3f",  x"0c", -- 0140
         x"3a",  x"07",  x"0d",  x"32",  x"3d",  x"0c",  x"cd",  x"70", -- 0148
         x"02",  x"cd",  x"f0",  x"05",  x"8a",  x"14",  x"cd",  x"f0", -- 0150
         x"05",  x"11",  x"15",  x"21",  x"b6",  x"f8",  x"22",  x"3f", -- 0158
         x"0c",  x"3a",  x"1a",  x"0d",  x"cd",  x"9b",  x"07",  x"3e", -- 0160
         x"1d",  x"fd",  x"cb",  x"00",  x"46",  x"20",  x"02",  x"3e", -- 0168
         x"15",  x"21",  x"c0",  x"f8",  x"cd",  x"bc",  x"01",  x"cd", -- 0170
         x"5a",  x"06",  x"2a",  x"01",  x"0d",  x"cd",  x"73",  x"06", -- 0178
         x"06",  x"0f",  x"2a",  x"01",  x"0d",  x"23",  x"36",  x"80", -- 0180
         x"10",  x"fb",  x"23",  x"36",  x"81",  x"06",  x"16",  x"23", -- 0188
         x"36",  x"91",  x"10",  x"fb",  x"04",  x"cd",  x"d1",  x"04", -- 0190
         x"cd",  x"73",  x"06",  x"06",  x"13",  x"fd",  x"cb",  x"00", -- 0198
         x"46",  x"20",  x"02",  x"06",  x"0b",  x"cd",  x"d1",  x"04", -- 01A0
         x"06",  x"01",  x"cd",  x"03",  x"06",  x"fd",  x"cb",  x"00", -- 01A8
         x"46",  x"28",  x"06",  x"21",  x"44",  x"15",  x"cd",  x"e0", -- 01B0
         x"01",  x"01",  x"2c",  x"01",  x"c5",  x"cd",  x"00",  x"04", -- 01B8
         x"3a",  x"bf",  x"0c",  x"b7",  x"20",  x"09",  x"3e",  x"4d", -- 01C0
         x"32",  x"bf",  x"0c",  x"21",  x"06",  x"0d",  x"34",  x"21", -- 01C8
         x"56",  x"0c",  x"3a",  x"05",  x"0d",  x"c6",  x"01",  x"38", -- 01D0
         x"0b",  x"fe",  x"02",  x"28",  x"07",  x"fe",  x"01",  x"20", -- 01D8
         x"09",  x"35",  x"28",  x"05",  x"35",  x"28",  x"02",  x"18", -- 01E0
         x"01",  x"34",  x"06",  x"08",  x"cd",  x"c7",  x"01",  x"10", -- 01E8
         x"fb",  x"fd",  x"cb",  x"00",  x"46",  x"ca",  x"8f",  x"13", -- 01F0
         x"21",  x"58",  x"0d",  x"3a",  x"56",  x"0c",  x"c6",  x"18", -- 01F8
         x"77",  x"2b",  x"cd",  x"d4",  x"01",  x"21",  x"20",  x"f8", -- 0200
         x"22",  x"3f",  x"0c",  x"3a",  x"06",  x"0d",  x"32",  x"3d", -- 0208
         x"0c",  x"cd",  x"70",  x"02",  x"36",  x"20",  x"2b",  x"36", -- 0210
         x"20",  x"2b",  x"36",  x"2c",  x"c1",  x"0b",  x"21",  x"3a", -- 0218
         x"f8",  x"22",  x"3f",  x"0c",  x"ed",  x"43",  x"3d",  x"0c", -- 0220
         x"cd",  x"70",  x"02",  x"78",  x"b1",  x"20",  x"8d",  x"3a", -- 0228
         x"bf",  x"0c",  x"47",  x"3a",  x"06",  x"0d",  x"dd",  x"77", -- 0230
         x"06",  x"3e",  x"50",  x"90",  x"dd",  x"77",  x"05",  x"32", -- 0238
         x"3d",  x"0c",  x"21",  x"22",  x"f8",  x"36",  x"2c",  x"23", -- 0240
         x"22",  x"3f",  x"0c",  x"cd",  x"70",  x"02",  x"36",  x"45", -- 0248
         x"2b",  x"36",  x"53",  x"21",  x"20",  x"f8",  x"7e",  x"dd", -- 0250
         x"77",  x"01",  x"23",  x"7e",  x"dd",  x"77",  x"02",  x"23", -- 0258
         x"23",  x"7e",  x"dd",  x"77",  x"03",  x"23",  x"7e",  x"dd", -- 0260
         x"77",  x"04",  x"fd",  x"cb",  x"00",  x"46",  x"28",  x"06", -- 0268
         x"21",  x"e1",  x"15",  x"cd",  x"d4",  x"01",  x"21",  x"1a", -- 0270
         x"0d",  x"7e",  x"dd",  x"77",  x"00",  x"cb",  x"2e",  x"3e", -- 0278
         x"01",  x"be",  x"38",  x"01",  x"77",  x"21",  x"c3",  x"fa", -- 0280
         x"11",  x"40",  x"00",  x"06",  x"03",  x"cd",  x"56",  x"07", -- 0288
         x"19",  x"10",  x"fa",  x"06",  x"04",  x"21",  x"92",  x"14", -- 0290
         x"c5",  x"cd",  x"f8",  x"05",  x"c1",  x"10",  x"f9",  x"21", -- 0298
         x"83",  x"fb",  x"11",  x"40",  x"00",  x"0e",  x"31",  x"dd", -- 02A0
         x"21",  x"1d",  x"0d",  x"3a",  x"07",  x"0d",  x"47",  x"cd", -- 02A8
         x"62",  x"07",  x"19",  x"cd",  x"62",  x"07",  x"e5",  x"d5", -- 02B0
         x"11",  x"04",  x"00",  x"19",  x"71",  x"0c",  x"11",  x"06", -- 02B8
         x"00",  x"19",  x"22",  x"3f",  x"0c",  x"dd",  x"7e",  x"00", -- 02C0
         x"cd",  x"9b",  x"07",  x"c5",  x"11",  x"06",  x"00",  x"19", -- 02C8
         x"dd",  x"7e",  x"01",  x"77",  x"23",  x"dd",  x"7e",  x"02", -- 02D0
         x"77",  x"23",  x"36",  x"2c",  x"23",  x"dd",  x"7e",  x"03", -- 02D8
         x"77",  x"23",  x"dd",  x"7e",  x"04",  x"77",  x"23",  x"11", -- 02E0
         x"24",  x"15",  x"cd",  x"90",  x"07",  x"11",  x"05",  x"00", -- 02E8
         x"19",  x"22",  x"3f",  x"0c",  x"dd",  x"6e",  x"05",  x"dd", -- 02F0
         x"66",  x"06",  x"7d",  x"b4",  x"20",  x"09",  x"2a",  x"3f", -- 02F8
         x"0c",  x"2b",  x"11",  x"36",  x"15",  x"18",  x"59",  x"cb", -- 0300
         x"25",  x"11",  x"00",  x"50",  x"eb",  x"ed",  x"52",  x"44", -- 0308
         x"0e",  x"00",  x"e5",  x"d1",  x"19",  x"30",  x"01",  x"0c", -- 0310
         x"10",  x"fa",  x"cb",  x"25",  x"cb",  x"14",  x"cb",  x"11", -- 0318
         x"cb",  x"25",  x"cb",  x"14",  x"cb",  x"11",  x"6c",  x"61", -- 0320
         x"dd",  x"5e",  x"00",  x"af",  x"57",  x"47",  x"4f",  x"ed", -- 0328
         x"52",  x"03",  x"30",  x"fb",  x"21",  x"e8",  x"03",  x"ed", -- 0330
         x"42",  x"38",  x"07",  x"2a",  x"3f",  x"0c",  x"23",  x"22", -- 0338
         x"3f",  x"0c",  x"ed",  x"43",  x"3d",  x"0c",  x"2a",  x"0e", -- 0340
         x"0c",  x"b7",  x"ed",  x"42",  x"30",  x"0a",  x"fd",  x"cb", -- 0348
         x"00",  x"46",  x"28",  x"04",  x"ed",  x"43",  x"0e",  x"0c", -- 0350
         x"cd",  x"70",  x"02",  x"2b",  x"2b",  x"11",  x"2e",  x"15", -- 0358
         x"cd",  x"90",  x"07",  x"01",  x"07",  x"00",  x"dd",  x"09", -- 0360
         x"c1",  x"d1",  x"e1",  x"19",  x"05",  x"c2",  x"af",  x"12", -- 0368
         x"cd",  x"62",  x"07",  x"19",  x"cd",  x"56",  x"07",  x"06", -- 0370
         x"03",  x"cd",  x"03",  x"06",  x"fd",  x"cb",  x"00",  x"46", -- 0378
         x"c2",  x"ef",  x"10",  x"21",  x"07",  x"0d",  x"7e",  x"fe", -- 0380
         x"03",  x"da",  x"ef",  x"10",  x"c3",  x"73",  x"10",  x"06", -- 0388
         x"60",  x"c5",  x"cd",  x"9a",  x"01",  x"c1",  x"c2",  x"f1", -- 0390
         x"00",  x"3a",  x"03",  x"0c",  x"b7",  x"c2",  x"00",  x"10", -- 0398
         x"10",  x"ef",  x"c3",  x"05",  x"12",  x"9b",  x"98",  x"95", -- 03A0
         x"92",  x"8f",  x"8c",  x"89",  x"86",  x"83",  x"00",  x"f8", -- 03A8
         x"3d",  x"3d",  x"3d",  x"20",  x"52",  x"45",  x"4b",  x"4f", -- 03B0
         x"52",  x"44",  x"3a",  x"20",  x"30",  x"30",  x"20",  x"3d", -- 03B8
         x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d", -- 03C0
         x"3d",  x"3d",  x"20",  x"5a",  x"45",  x"49",  x"54",  x"3a", -- 03C8
         x"20",  x"30",  x"30",  x"2c",  x"30",  x"30",  x"20",  x"53", -- 03D0
         x"45",  x"4b",  x"2e",  x"20",  x"3d",  x"3d",  x"3d",  x"20", -- 03D8
         x"45",  x"4e",  x"54",  x"46",  x"2e",  x"5a",  x"49",  x"45", -- 03E0
         x"4c",  x"3a",  x"20",  x"3d",  x"3d",  x"3d",  x"10",  x"fc", -- 03E8
         x"2f",  x"57",  x"55",  x"45",  x"4e",  x"53",  x"43",  x"48", -- 03F0
         x"45",  x"4e",  x"20",  x"53",  x"49",  x"45",  x"20",  x"45"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
