library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom2_4000 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom2_4000;

architecture rtl of rom2_4000 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"3e",  x"79",  x"32",  x"38",  x"0d",  x"3e",  x"4d",  x"32", -- 0000
         x"bf",  x"0c",  x"fd",  x"21",  x"36",  x"0d",  x"fd",  x"36", -- 0008
         x"01",  x"0f",  x"cd",  x"b7",  x"02",  x"21",  x"71",  x"48", -- 0010
         x"11",  x"10",  x"f4",  x"ed",  x"4b",  x"f0",  x"4a",  x"ed", -- 0018
         x"b0",  x"21",  x"f2",  x"4a",  x"11",  x"00",  x"f0",  x"ed", -- 0020
         x"4b",  x"ea",  x"4d",  x"ed",  x"b0",  x"21",  x"ec",  x"4d", -- 0028
         x"11",  x"30",  x"ec",  x"ed",  x"4b",  x"8c",  x"4e",  x"ed", -- 0030
         x"b0",  x"21",  x"8e",  x"4e",  x"11",  x"10",  x"ed",  x"ed", -- 0038
         x"4b",  x"ea",  x"4f",  x"ed",  x"b0",  x"21",  x"00",  x"f8", -- 0040
         x"11",  x"01",  x"f8",  x"36",  x"81",  x"01",  x"ff",  x"07", -- 0048
         x"ed",  x"b0",  x"cd",  x"74",  x"44",  x"ff",  x"46",  x"01", -- 0050
         x"0e",  x"00",  x"62",  x"6b",  x"36",  x"ce",  x"13",  x"ed", -- 0058
         x"b0",  x"21",  x"bd",  x"ff",  x"22",  x"3c",  x"0d",  x"36", -- 0060
         x"de",  x"23",  x"36",  x"de",  x"2a",  x"0a",  x"0c",  x"22", -- 0068
         x"3d",  x"0c",  x"21",  x"0a",  x"f8",  x"22",  x"3f",  x"0c", -- 0070
         x"cd",  x"70",  x"02",  x"3e",  x"82",  x"dd",  x"21",  x"a1", -- 0078
         x"47",  x"06",  x"03",  x"c5",  x"06",  x"06",  x"cd",  x"d0", -- 0080
         x"42",  x"10",  x"fb",  x"c1",  x"c6",  x"04",  x"10",  x"f3", -- 0088
         x"dd",  x"21",  x"c5",  x"47",  x"dd",  x"6e",  x"00",  x"dd", -- 0090
         x"66",  x"01",  x"22",  x"32",  x"0d",  x"af",  x"32",  x"34", -- 0098
         x"0d",  x"3e",  x"02",  x"32",  x"35",  x"0d",  x"dd",  x"21", -- 00A0
         x"32",  x"0d",  x"3e",  x"b6",  x"cd",  x"f0",  x"42",  x"01", -- 00A8
         x"0f",  x"05",  x"21",  x"cf",  x"47",  x"11",  x"00",  x"0d", -- 00B0
         x"ed",  x"a0",  x"ed",  x"a0",  x"cd",  x"4a",  x"44",  x"10", -- 00B8
         x"f7",  x"11",  x"08",  x"00",  x"dd",  x"21",  x"00",  x"0d", -- 00C0
         x"06",  x"05",  x"dd",  x"7e",  x"02",  x"cd",  x"d0",  x"42", -- 00C8
         x"dd",  x"19",  x"10",  x"f6",  x"dd",  x"21",  x"00",  x"0d", -- 00D0
         x"06",  x"05",  x"e5",  x"2a",  x"18",  x"0c",  x"22",  x"3d", -- 00D8
         x"0c",  x"21",  x"1a",  x"f8",  x"22",  x"3f",  x"0c",  x"cd", -- 00E0
         x"70",  x"02",  x"e1",  x"af",  x"c5",  x"dd",  x"be",  x"05", -- 00E8
         x"c2",  x"5c",  x"41",  x"dd",  x"35",  x"03",  x"fa",  x"64", -- 00F0
         x"41",  x"3e",  x"03",  x"dd",  x"be",  x"03",  x"c2",  x"5f", -- 00F8
         x"41",  x"ed",  x"5f",  x"e6",  x"0e",  x"21",  x"d9",  x"47", -- 0100
         x"85",  x"6f",  x"30",  x"01",  x"24",  x"5e",  x"23",  x"56", -- 0108
         x"eb",  x"dd",  x"5e",  x"00",  x"dd",  x"56",  x"01",  x"dd", -- 0110
         x"cb",  x"04",  x"46",  x"28",  x"16",  x"6b",  x"62",  x"dd", -- 0118
         x"35",  x"04",  x"06",  x"81",  x"cd",  x"a7",  x"43",  x"38", -- 0120
         x"2e",  x"06",  x"92",  x"cd",  x"a7",  x"43",  x"c2",  x"8f", -- 0128
         x"41",  x"18",  x"24",  x"19",  x"cd",  x"ad",  x"42",  x"06", -- 0130
         x"81",  x"cd",  x"a7",  x"43",  x"38",  x"19",  x"06",  x"92", -- 0138
         x"cd",  x"a7",  x"43",  x"28",  x"4a",  x"fe",  x"82",  x"28", -- 0140
         x"23",  x"fe",  x"86",  x"28",  x"1f",  x"fe",  x"8a",  x"28", -- 0148
         x"1b",  x"fe",  x"8e",  x"28",  x"17",  x"18",  x"1c",  x"cd", -- 0150
         x"d3",  x"46",  x"18",  x"03",  x"dd",  x"35",  x"05",  x"11", -- 0158
         x"0a",  x"00",  x"18",  x"34",  x"3e",  x"92",  x"dd",  x"36", -- 0160
         x"03",  x"05",  x"18",  x"26",  x"ed",  x"5f",  x"c6",  x"40", -- 0168
         x"dd",  x"77",  x"05",  x"dd",  x"75",  x"00",  x"dd",  x"74", -- 0170
         x"01",  x"7e",  x"dd",  x"77",  x"06",  x"23",  x"7e",  x"dd", -- 0178
         x"77",  x"07",  x"11",  x"3f",  x"00",  x"19",  x"7e",  x"dd", -- 0180
         x"77",  x"08",  x"23",  x"7e",  x"dd",  x"77",  x"09",  x"dd", -- 0188
         x"7e",  x"02",  x"cd",  x"d0",  x"42",  x"11",  x"08",  x"00", -- 0190
         x"dd",  x"19",  x"c1",  x"05",  x"c2",  x"eb",  x"40",  x"fd", -- 0198
         x"cb",  x"01",  x"4e",  x"c2",  x"1f",  x"42",  x"db",  x"84", -- 01A0
         x"fd",  x"77",  x"00",  x"dd",  x"21",  x"32",  x"0d",  x"dd", -- 01A8
         x"35",  x"03",  x"20",  x"2d",  x"dd",  x"36",  x"03",  x"02", -- 01B0
         x"dd",  x"5e",  x"00",  x"dd",  x"56",  x"01",  x"fd",  x"cb", -- 01B8
         x"00",  x"1e",  x"cd",  x"ed",  x"44",  x"fd",  x"cb",  x"00", -- 01C0
         x"1e",  x"d4",  x"54",  x"46",  x"fd",  x"cb",  x"00",  x"1e", -- 01C8
         x"d4",  x"b2",  x"46",  x"fd",  x"cb",  x"00",  x"1e",  x"d4", -- 01D0
         x"c9",  x"46",  x"fd",  x"cb",  x"00",  x"1e",  x"d4",  x"ce", -- 01D8
         x"46",  x"cd",  x"87",  x"44",  x"c2",  x"d4",  x"40",  x"af", -- 01E0
         x"32",  x"03",  x"0c",  x"21",  x"80",  x"fb",  x"36",  x"20", -- 01E8
         x"54",  x"5d",  x"13",  x"01",  x"3f",  x"01",  x"ed",  x"b0", -- 01F0
         x"2a",  x"18",  x"0c",  x"ed",  x"5b",  x"0a",  x"0c",  x"b7", -- 01F8
         x"ed",  x"52",  x"38",  x"14",  x"cd",  x"74",  x"44",  x"3f", -- 0200
         x"47",  x"2a",  x"18",  x"0c",  x"22",  x"0a",  x"0c",  x"21", -- 0208
         x"f6",  x"47",  x"cd",  x"e0",  x"01",  x"c3",  x"f1",  x"00", -- 0210
         x"cd",  x"74",  x"44",  x"33",  x"47",  x"18",  x"f0",  x"fd", -- 0218
         x"cb",  x"01",  x"7e",  x"20",  x"57",  x"fd",  x"36",  x"01", -- 0220
         x"ff",  x"21",  x"00",  x"fc",  x"3e",  x"10",  x"cd",  x"bc", -- 0228
         x"01",  x"cd",  x"74",  x"44",  x"4e",  x"47",  x"11",  x"92", -- 0230
         x"ff",  x"21",  x"0a",  x"03",  x"01",  x"1b",  x"00",  x"ed", -- 0238
         x"b0",  x"21",  x"44",  x"fd",  x"06",  x"04",  x"11",  x"59", -- 0240
         x"48",  x"c5",  x"0e",  x"04",  x"1a",  x"13",  x"47",  x"36", -- 0248
         x"81",  x"23",  x"10",  x"fb",  x"1a",  x"13",  x"85",  x"6f", -- 0250
         x"30",  x"01",  x"24",  x"0d",  x"20",  x"ee",  x"c1",  x"10", -- 0258
         x"e5",  x"dd",  x"21",  x"61",  x"48",  x"06",  x"08",  x"3e", -- 0260
         x"96",  x"cd",  x"d0",  x"42",  x"c6",  x"04",  x"10",  x"f9", -- 0268
         x"06",  x"04",  x"21",  x"66",  x"47",  x"c5",  x"cd",  x"7c", -- 0270
         x"44",  x"c1",  x"10",  x"f9",  x"cd",  x"c7",  x"01",  x"cd", -- 0278
         x"c7",  x"01",  x"af",  x"32",  x"56",  x"0c",  x"cd",  x"9a", -- 0280
         x"01",  x"c2",  x"f1",  x"00",  x"3a",  x"03",  x"0c",  x"b7", -- 0288
         x"ca",  x"d4",  x"40",  x"fd",  x"36",  x"01",  x"00",  x"21", -- 0290
         x"38",  x"48",  x"cd",  x"e0",  x"01",  x"2a",  x"00",  x"0c", -- 0298
         x"23",  x"22",  x"00",  x"0c",  x"21",  x"00",  x"00",  x"22", -- 02A0
         x"18",  x"0c",  x"c3",  x"45",  x"40",  x"f5",  x"d5",  x"e5", -- 02A8
         x"dd",  x"6e",  x"00",  x"dd",  x"66",  x"01",  x"11",  x"3f", -- 02B0
         x"00",  x"dd",  x"7e",  x"06",  x"77",  x"23",  x"dd",  x"7e", -- 02B8
         x"07",  x"77",  x"19",  x"dd",  x"7e",  x"08",  x"77",  x"23", -- 02C0
         x"dd",  x"7e",  x"09",  x"77",  x"e1",  x"d1",  x"f1",  x"c9", -- 02C8
         x"d5",  x"f5",  x"e5",  x"c5",  x"01",  x"3f",  x"00",  x"dd", -- 02D0
         x"6e",  x"00",  x"dd",  x"66",  x"01",  x"dd",  x"23",  x"dd", -- 02D8
         x"23",  x"77",  x"3c",  x"23",  x"77",  x"3c",  x"09",  x"77", -- 02E0
         x"3c",  x"23",  x"77",  x"c1",  x"e1",  x"f1",  x"d1",  x"c9", -- 02E8
         x"d5",  x"16",  x"01",  x"cd",  x"8e",  x"43",  x"f5",  x"1e", -- 02F0
         x"04",  x"e5",  x"c5",  x"01",  x"3e",  x"00",  x"dd",  x"6e", -- 02F8
         x"00",  x"dd",  x"66",  x"01",  x"77",  x"82",  x"23",  x"77", -- 0300
         x"82",  x"23",  x"77",  x"82",  x"09",  x"1d",  x"20",  x"f4", -- 0308
         x"18",  x"d9",  x"d5",  x"16",  x"00",  x"cd",  x"1a",  x"43", -- 0310
         x"18",  x"dc",  x"d5",  x"f5",  x"16",  x"00",  x"e5",  x"c5", -- 0318
         x"01",  x"c0",  x"ff",  x"dd",  x"6e",  x"00",  x"dd",  x"66", -- 0320
         x"01",  x"09",  x"dd",  x"cb",  x"02",  x"5e",  x"20",  x"68", -- 0328
         x"2b",  x"2b",  x"01",  x"01",  x"00",  x"cb",  x"42",  x"28", -- 0330
         x"3d",  x"3e",  x"d2",  x"5e",  x"dd",  x"e5",  x"dd",  x"21", -- 0338
         x"46",  x"0d",  x"cd",  x"67",  x"43",  x"dd",  x"73",  x"00", -- 0340
         x"77",  x"09",  x"82",  x"5e",  x"cd",  x"67",  x"43",  x"dd", -- 0348
         x"73",  x"01",  x"77",  x"01",  x"40",  x"00",  x"09",  x"82", -- 0350
         x"5e",  x"cd",  x"67",  x"43",  x"dd",  x"73",  x"02",  x"dd", -- 0358
         x"e1",  x"77",  x"c1",  x"e1",  x"f1",  x"d1",  x"c9",  x"f5", -- 0360
         x"3e",  x"91",  x"bb",  x"38",  x"02",  x"f1",  x"c9",  x"f1", -- 0368
         x"e3",  x"23",  x"23",  x"23",  x"e3",  x"c9",  x"dd",  x"e5", -- 0370
         x"dd",  x"21",  x"46",  x"0d",  x"dd",  x"7e",  x"00",  x"77", -- 0378
         x"09",  x"dd",  x"7e",  x"01",  x"77",  x"01",  x"40",  x"00", -- 0380
         x"09",  x"dd",  x"7e",  x"02",  x"18",  x"d1",  x"d5",  x"f5", -- 0388
         x"16",  x"01",  x"af",  x"32",  x"39",  x"0d",  x"18",  x"86", -- 0390
         x"01",  x"04",  x"00",  x"09",  x"01",  x"ff",  x"ff",  x"cb", -- 0398
         x"42",  x"28",  x"d3",  x"3e",  x"d8",  x"18",  x"94",  x"e5", -- 03A0
         x"d5",  x"c5",  x"0e",  x"00",  x"7e",  x"cd",  x"c9",  x"43", -- 03A8
         x"23",  x"7e",  x"cd",  x"c9",  x"43",  x"11",  x"3f",  x"00", -- 03B0
         x"19",  x"7e",  x"cd",  x"c9",  x"43",  x"23",  x"7e",  x"cd", -- 03B8
         x"c9",  x"43",  x"c5",  x"f1",  x"c1",  x"d1",  x"e1",  x"7e", -- 03C0
         x"c9",  x"b8",  x"38",  x"05",  x"79",  x"f6",  x"40",  x"4f", -- 03C8
         x"c9",  x"79",  x"f6",  x"01",  x"4f",  x"c9",  x"e5",  x"d5", -- 03D0
         x"c5",  x"0e",  x"00",  x"16",  x"04",  x"7d",  x"cd",  x"0f", -- 03D8
         x"44",  x"c6",  x"ff",  x"e6",  x"3f",  x"20",  x"02",  x"0e", -- 03E0
         x"01",  x"7e",  x"cd",  x"c9",  x"43",  x"23",  x"7e",  x"cd", -- 03E8
         x"c9",  x"43",  x"23",  x"7e",  x"cd",  x"c9",  x"43",  x"15", -- 03F0
         x"28",  x"08",  x"d5",  x"11",  x"3e",  x"00",  x"19",  x"d1"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
