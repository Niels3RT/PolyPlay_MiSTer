library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom2_2400 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom2_2400;

architecture rtl of rom2_2400 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"50",  x"12",  x"82",  x"01",  x"20",  x"dc",  x"82",  x"01", -- 0000
         x"08",  x"dc",  x"82",  x"01",  x"08",  x"c4",  x"82",  x"01", -- 0008
         x"08",  x"af",  x"82",  x"01",  x"08",  x"a5",  x"82",  x"01", -- 0010
         x"20",  x"93",  x"82",  x"01",  x"10",  x"af",  x"82",  x"01", -- 0018
         x"10",  x"af",  x"82",  x"01",  x"10",  x"c4",  x"82",  x"01", -- 0020
         x"10",  x"93",  x"82",  x"01",  x"10",  x"c4",  x"82",  x"01", -- 0028
         x"10",  x"93",  x"82",  x"01",  x"10",  x"af",  x"82",  x"01", -- 0030
         x"10",  x"c4",  x"82",  x"01",  x"10",  x"dc",  x"00",  x"00", -- 0038
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"10", -- 0040
         x"93",  x"82",  x"01",  x"10",  x"6b",  x"82",  x"01",  x"10", -- 0048
         x"93",  x"82",  x"01",  x"10",  x"93",  x"82",  x"01",  x"10", -- 0050
         x"af",  x"82",  x"01",  x"10",  x"af",  x"82",  x"01",  x"10", -- 0058
         x"c4",  x"82",  x"01",  x"20",  x"c4",  x"00",  x"20",  x"20", -- 0060
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0068
         x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0070
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0078
         x"ff",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0080
         x"00",  x"b5",  x"4a",  x"2d",  x"12",  x"1f",  x"04",  x"03", -- 0088
         x"01",  x"50",  x"a8",  x"48",  x"b0",  x"c0",  x"80",  x"e0", -- 0090
         x"fe",  x"00",  x"00",  x"00",  x"3f",  x"ff",  x"ff",  x"ff", -- 0098
         x"ff",  x"00",  x"00",  x"01",  x"ff",  x"ff",  x"ff",  x"ff", -- 00A0
         x"ff",  x"df",  x"fe",  x"fc",  x"f0",  x"f0",  x"f0",  x"f0", -- 00A8
         x"e0",  x"7f",  x"7f",  x"30",  x"50",  x"50",  x"90",  x"90", -- 00B0
         x"90",  x"ff",  x"ff",  x"03",  x"03",  x"02",  x"02",  x"02", -- 00B8
         x"02",  x"c0",  x"80",  x"00",  x"00",  x"80",  x"40",  x"20", -- 00C0
         x"20",  x"7f",  x"7f",  x"30",  x"28",  x"28",  x"24",  x"24", -- 00C8
         x"28",  x"ff",  x"ff",  x"03",  x"03",  x"05",  x"05",  x"09", -- 00D0
         x"11",  x"c0",  x"80",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00D8
         x"00",  x"0a",  x"15",  x"12",  x"0d",  x"03",  x"01",  x"07", -- 00E0
         x"7f",  x"ad",  x"52",  x"b4",  x"48",  x"f8",  x"20",  x"c0", -- 00E8
         x"80",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00F0
         x"00",  x"fb",  x"7f",  x"3f",  x"0f",  x"0f",  x"0f",  x"0f", -- 00F8
         x"07",  x"00",  x"00",  x"80",  x"ff",  x"ff",  x"ff",  x"ff", -- 0100
         x"ff",  x"00",  x"00",  x"00",  x"fc",  x"ff",  x"ff",  x"ff", -- 0108
         x"ff",  x"03",  x"01",  x"00",  x"00",  x"01",  x"02",  x"04", -- 0110
         x"04",  x"ff",  x"ff",  x"c0",  x"c0",  x"40",  x"40",  x"40", -- 0118
         x"40",  x"fe",  x"fe",  x"0c",  x"0a",  x"0a",  x"09",  x"09", -- 0120
         x"09",  x"03",  x"01",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0128
         x"00",  x"ff",  x"ff",  x"c0",  x"c0",  x"a0",  x"a0",  x"90", -- 0130
         x"88",  x"fe",  x"fe",  x"0c",  x"14",  x"14",  x"24",  x"24", -- 0138
         x"14",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0140
         x"00",  x"00",  x"18",  x"18",  x"18",  x"18",  x"18",  x"18", -- 0148
         x"3c",  x"00",  x"00",  x"f4",  x"fc",  x"78",  x"30",  x"01", -- 0150
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"02",  x"ff", -- 0158
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0160
         x"ee",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0168
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"40",  x"ff", -- 0170
         x"00",  x"00",  x"00",  x"2f",  x"3f",  x"1e",  x"0c",  x"80", -- 0178
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0180
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0188
         x"77",  x"00",  x"00",  x"00",  x"00",  x"00",  x"06",  x"06", -- 0190
         x"00",  x"00",  x"01",  x"02",  x"01",  x"00",  x"00",  x"00", -- 0198
         x"3f",  x"25",  x"5a",  x"95",  x"67",  x"9c",  x"60",  x"01", -- 01A0
         x"ff",  x"40",  x"b0",  x"60",  x"fe",  x"df",  x"fe",  x"fc", -- 01A8
         x"f0",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f",  x"7f",  x"0e", -- 01B0
         x"fe",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"01", -- 01B8
         x"1f",  x"f0",  x"f0",  x"f0",  x"e0",  x"c0",  x"80",  x"80", -- 01C0
         x"80",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 01C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 01D0
         x"ff",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01E0
         x"00",  x"b5",  x"4a",  x"2d",  x"12",  x"1f",  x"04",  x"00", -- 01E8
         x"00",  x"50",  x"a8",  x"48",  x"b0",  x"c0",  x"80",  x"00", -- 01F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0200
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0208
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0210
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0218
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0220
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0228
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0230
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0238
         x"00",  x"0a",  x"15",  x"12",  x"0d",  x"03",  x"01",  x"00", -- 0240
         x"00",  x"ad",  x"52",  x"b4",  x"48",  x"f8",  x"20",  x"00", -- 0248
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0250
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0258
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0260
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0268
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0270
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0278
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0280
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0288
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0290
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0298
         x"00",  x"18",  x"3c",  x"3c",  x"7e",  x"7e",  x"ff",  x"ff", -- 02A0
         x"ff",  x"ff",  x"66",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02A8
         x"00",  x"78",  x"fe",  x"f4",  x"fc",  x"78",  x"30",  x"7e", -- 02B0
         x"fe",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02B8
         x"60",  x"ff",  x"fc",  x"78",  x"fc",  x"fc",  x"cc",  x"cc", -- 02C0
         x"00",  x"c0",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02D0
         x"06",  x"1e",  x"7f",  x"2f",  x"3f",  x"1e",  x"0c",  x"7e", -- 02D8
         x"7f",  x"03",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02E0
         x"00",  x"ff",  x"3f",  x"1e",  x"3f",  x"3f",  x"33",  x"33", -- 02E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"06",  x"06", -- 02F0
         x"00",  x"00",  x"01",  x"02",  x"01",  x"00",  x"00",  x"00", -- 02F8
         x"00",  x"25",  x"5a",  x"95",  x"60",  x"90",  x"60",  x"00", -- 0300
         x"00",  x"40",  x"b0",  x"60",  x"20",  x"04",  x"00",  x"00", -- 0308
         x"08",  x"00",  x"00",  x"10",  x"00",  x"00",  x"00",  x"00", -- 0310
         x"00",  x"06",  x"06",  x"00",  x"82",  x"3d",  x"0c",  x"81", -- 0318
         x"cd",  x"82",  x"70",  x"02",  x"81",  x"21",  x"82",  x"2b", -- 0320
         x"f8",  x"81",  x"22",  x"82",  x"3f",  x"0c",  x"81",  x"2a", -- 0328
         x"82",  x"1a",  x"0c",  x"81",  x"22",  x"82",  x"3d",  x"0c", -- 0330
         x"81",  x"cd",  x"82",  x"70",  x"02",  x"81",  x"21",  x"82", -- 0338
         x"3b",  x"f8",  x"81",  x"22",  x"82",  x"3f",  x"0c",  x"81", -- 0340
         x"3a",  x"82",  x"e4",  x"0c",  x"81",  x"26",  x"81",  x"00", -- 0348
         x"81",  x"6f",  x"81",  x"22",  x"82",  x"3d",  x"0c",  x"81", -- 0350
         x"cd",  x"82",  x"70",  x"02",  x"81",  x"c9",  x"81",  x"e5", -- 0358
         x"81",  x"2a",  x"82",  x"cb",  x"0c",  x"81",  x"cd",  x"82", -- 0360
         x"b5",  x"32",  x"81",  x"ed",  x"81",  x"43",  x"82",  x"ce", -- 0368
         x"0c",  x"81",  x"e1",  x"81",  x"c9",  x"81",  x"e5",  x"81", -- 0370
         x"5e",  x"81",  x"23",  x"81",  x"56",  x"81",  x"eb",  x"81", -- 0378
         x"cd",  x"82",  x"b5",  x"32",  x"81",  x"e1",  x"81",  x"23", -- 0380
         x"81",  x"23",  x"81",  x"71",  x"81",  x"23",  x"81",  x"70", -- 0388
         x"81",  x"2b",  x"81",  x"2b",  x"81",  x"2b",  x"81",  x"c9", -- 0390
         x"81",  x"11",  x"82",  x"00",  x"f8",  x"81",  x"01",  x"82", -- 0398
         x"00",  x"00",  x"81",  x"af",  x"81",  x"ed",  x"81",  x"52", -- 03A0
         x"81",  x"11",  x"82",  x"40",  x"00",  x"81",  x"af",  x"81", -- 03A8
         x"ed",  x"81",  x"52",  x"81",  x"c8",  x"81",  x"38",  x"81", -- 03B0
         x"03",  x"81",  x"04",  x"81",  x"18",  x"81",  x"f7",  x"81", -- 03B8
         x"ed",  x"81",  x"5a",  x"81",  x"4d",  x"81",  x"c9",  x"81", -- 03C0
         x"2a",  x"82",  x"93",  x"0c",  x"81",  x"23",  x"81",  x"23", -- 03C8
         x"81",  x"4e",  x"81",  x"23",  x"81",  x"46",  x"81",  x"21", -- 03D0
         x"82",  x"00",  x"f8",  x"81",  x"11",  x"82",  x"40",  x"00", -- 03D8
         x"81",  x"af",  x"81",  x"b8",  x"81",  x"28",  x"81",  x"05", -- 03E0
         x"81",  x"05",  x"81",  x"19",  x"81",  x"d8",  x"81",  x"18", -- 03E8
         x"81",  x"f7",  x"81",  x"09",  x"81",  x"2b",  x"81",  x"eb", -- 03F0
         x"81",  x"2a",  x"82",  x"93",  x"0c",  x"81",  x"73",  x"81"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
