library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom2_1800 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom2_1800;

architecture rtl of rom2_1800 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"00",  x"00",  x"00",  x"00",  x"00",  x"18",  x"18",  x"00", -- 0000
         x"00",  x"00",  x"d8",  x"00",  x"01",  x"00",  x"00",  x"3c", -- 0008
         x"7e",  x"7e",  x"7e",  x"3c",  x"00",  x"10",  x"00",  x"07", -- 0010
         x"18",  x"00",  x"7e",  x"5a",  x"66",  x"3c",  x"81",  x"42", -- 0018
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0020
         x"00",  x"00",  x"00",  x"00",  x"01",  x"00",  x"01",  x"00", -- 0028
         x"ff",  x"cb",  x"c3",  x"ff",  x"00",  x"00",  x"ff",  x"00", -- 0030
         x"00",  x"00",  x"00",  x"00",  x"80",  x"00",  x"80",  x"00", -- 0038
         x"03",  x"07",  x"01",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0040
         x"00",  x"c0",  x"e0",  x"c0",  x"00",  x"00",  x"00",  x"00", -- 0048
         x"28",  x"00",  x"05",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0050
         x"03",  x"cc",  x"33",  x"00",  x"03",  x"0c",  x"33",  x"cc", -- 0058
         x"30",  x"c0",  x"00",  x"cc",  x"30",  x"c0",  x"00",  x"00", -- 0060
         x"00",  x"00",  x"00",  x"03",  x"07",  x"01",  x"00",  x"00", -- 0068
         x"00",  x"00",  x"00",  x"00",  x"c0",  x"e0",  x"80",  x"00", -- 0070
         x"00",  x"00",  x"00",  x"10",  x"00",  x"08",  x"00",  x"00", -- 0078
         x"00",  x"00",  x"00",  x"00",  x"01",  x"03",  x"00",  x"00", -- 0080
         x"00",  x"00",  x"66",  x"cc",  x"b0",  x"60",  x"00",  x"00", -- 0088
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0090
         x"00",  x"00",  x"00",  x"00",  x"01",  x"0f",  x"06",  x"0d", -- 0098
         x"1b",  x"36",  x"6c",  x"d8",  x"b0",  x"60",  x"c0",  x"80", -- 00A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"03", -- 00A8
         x"07",  x"03",  x"00",  x"00",  x"00",  x"00",  x"00",  x"c0", -- 00B0
         x"e0",  x"c0",  x"00",  x"00",  x"00",  x"00",  x"30",  x"00", -- 00B8
         x"07",  x"00",  x"00",  x"66",  x"66",  x"66",  x"66",  x"66", -- 00C0
         x"66",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00C8
         x"00",  x"00",  x"03",  x"07",  x"03",  x"00",  x"00",  x"00", -- 00D0
         x"00",  x"c0",  x"e0",  x"c0",  x"00",  x"00",  x"00",  x"00", -- 00D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"36",  x"1b",  x"0d", -- 00E8
         x"06",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"80", -- 00F0
         x"c0",  x"10",  x"00",  x"07",  x"03",  x"01",  x"00",  x"00", -- 00F8
         x"00",  x"00",  x"00",  x"00",  x"60",  x"b0",  x"d8",  x"6c", -- 0100
         x"36",  x"1b",  x"0d",  x"06",  x"00",  x"00",  x"00",  x"00", -- 0108
         x"00",  x"00",  x"80",  x"f0",  x"00",  x"03",  x"07",  x"03", -- 0110
         x"00",  x"00",  x"00",  x"00",  x"c0",  x"e0",  x"c0",  x"00", -- 0118
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0120
         x"00",  x"00",  x"01",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0128
         x"00",  x"00",  x"80",  x"cc",  x"18",  x"00",  x"0b",  x"33", -- 0130
         x"0c",  x"03",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0138
         x"c0",  x"30",  x"cc",  x"33",  x"0c",  x"03",  x"00",  x"00", -- 0140
         x"00",  x"00",  x"00",  x"00",  x"c0",  x"33",  x"cc",  x"00", -- 0148
         x"00",  x"1f",  x"3f",  x"7f",  x"ff",  x"88",  x"ff",  x"01", -- 0150
         x"03",  x"ff",  x"7f",  x"7e",  x"7e",  x"70",  x"f0",  x"80", -- 0158
         x"c0",  x"ff",  x"fe",  x"3e",  x"3e",  x"06",  x"07",  x"00", -- 0160
         x"00",  x"f8",  x"fc",  x"fe",  x"ff",  x"11",  x"ff",  x"ff", -- 0168
         x"ff",  x"fc",  x"f8",  x"01",  x"01",  x"00",  x"00",  x"fe", -- 0170
         x"fe",  x"3f",  x"1f",  x"80",  x"80",  x"00",  x"00",  x"3f", -- 0178
         x"3f",  x"fc",  x"f8",  x"01",  x"01",  x"00",  x"00",  x"ff", -- 0180
         x"ff",  x"3f",  x"1f",  x"80",  x"80",  x"00",  x"00",  x"10", -- 0188
         x"01",  x"01",  x"18",  x"3c",  x"7e",  x"ff",  x"ff",  x"7e", -- 0190
         x"3c",  x"18",  x"d8",  x"00",  x"42",  x"00",  x"00",  x"3c", -- 0198
         x"7e",  x"7e",  x"7e",  x"3c",  x"00",  x"00",  x"00",  x"00", -- 01A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01A8
         x"00",  x"00",  x"00",  x"03",  x"07",  x"00",  x"00",  x"00", -- 01B0
         x"5a",  x"7e",  x"3c",  x"ff",  x"ff",  x"00",  x"00",  x"00", -- 01B8
         x"00",  x"00",  x"00",  x"c0",  x"e0",  x"07",  x"cd",  x"79", -- 01C0
         x"31",  x"01",  x"01",  x"00",  x"01",  x"ff",  x"cb",  x"c3", -- 01C8
         x"ff",  x"ff",  x"ff",  x"00",  x"ff",  x"e0",  x"b3",  x"be", -- 01D0
         x"9c",  x"80",  x"80",  x"00",  x"80",  x"03",  x"07",  x"03", -- 01D8
         x"02",  x"04",  x"04",  x"08",  x"08",  x"00",  x"c0",  x"e0", -- 01E0
         x"c0",  x"40",  x"40",  x"80",  x"80",  x"10",  x"10",  x"20", -- 01E8
         x"20",  x"40",  x"40",  x"f0",  x"40",  x"01",  x"03",  x"07", -- 01F0
         x"0f",  x"1e",  x"1e",  x"0e",  x"07",  x"ff",  x"fe",  x"bc", -- 01F8
         x"78",  x"78",  x"f0",  x"70",  x"38",  x"00",  x"01",  x"01", -- 0200
         x"01",  x"02",  x"02",  x"02",  x"07",  x"80",  x"00",  x"00", -- 0208
         x"00",  x"00",  x"00",  x"00",  x"c0",  x"03",  x"01",  x"00", -- 0210
         x"00",  x"01",  x"03",  x"cc",  x"33",  x"38",  x"9f",  x"fe", -- 0218
         x"ff",  x"dc",  x"30",  x"c0",  x"00",  x"cd",  x"30",  x"c0", -- 0220
         x"00",  x"00",  x"00",  x"00",  x"00",  x"03",  x"07",  x"03", -- 0228
         x"02",  x"02",  x"02",  x"04",  x"04",  x"00",  x"c0",  x"e0", -- 0230
         x"c0",  x"40",  x"40",  x"40",  x"80",  x"04",  x"04",  x"08", -- 0238
         x"08",  x"08",  x"08",  x"3e",  x"08",  x"01",  x"03",  x"07", -- 0240
         x"0f",  x"1e",  x"1e",  x"07",  x"03",  x"ff",  x"fe",  x"bc", -- 0248
         x"78",  x"78",  x"f0",  x"39",  x"9f",  x"00",  x"00",  x"00", -- 0250
         x"00",  x"66",  x"cc",  x"b0",  x"63",  x"80",  x"80",  x"80", -- 0258
         x"80",  x"80",  x"80",  x"80",  x"c0",  x"00",  x"00",  x"00", -- 0260
         x"00",  x"00",  x"00",  x"01",  x"0f",  x"ce",  x"6d",  x"3b", -- 0268
         x"36",  x"6c",  x"d8",  x"b0",  x"60",  x"c1",  x"81",  x"00", -- 0270
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"03",  x"07", -- 0278
         x"03",  x"01",  x"01",  x"01",  x"01",  x"00",  x"c0",  x"e0", -- 0280
         x"c0",  x"80",  x"80",  x"80",  x"80",  x"01",  x"01",  x"01", -- 0288
         x"01",  x"01",  x"01",  x"07",  x"01",  x"01",  x"01",  x"00", -- 0290
         x"00",  x"00",  x"00",  x"c0",  x"00",  x"ff",  x"e7",  x"e7", -- 0298
         x"e7",  x"e7",  x"e7",  x"e7",  x"e7",  x"80",  x"80",  x"00", -- 02A0
         x"00",  x"00",  x"00",  x"03",  x"00",  x"80",  x"80",  x"80", -- 02A8
         x"80",  x"80",  x"80",  x"e0",  x"80",  x"00",  x"00",  x"00", -- 02B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"e7",  x"e7",  x"e7", -- 02B8
         x"66",  x"66",  x"66",  x"66",  x"42",  x"00",  x"00",  x"00", -- 02C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"03",  x"07", -- 02C8
         x"03",  x"01",  x"01",  x"01",  x"01",  x"c0",  x"e0",  x"c0", -- 02D0
         x"40",  x"40",  x"40",  x"20",  x"20",  x"02",  x"02",  x"02", -- 02D8
         x"02",  x"02",  x"02",  x"0f",  x"04",  x"00",  x"00",  x"00", -- 02E0
         x"00",  x"36",  x"1b",  x"0d",  x"06",  x"ff",  x"7f",  x"3d", -- 02E8
         x"1e",  x"1e",  x"0f",  x"9c",  x"f9",  x"80",  x"c0",  x"e0", -- 02F0
         x"f0",  x"78",  x"78",  x"e0",  x"c0",  x"20",  x"20",  x"20", -- 02F8
         x"10",  x"10",  x"10",  x"7c",  x"10",  x"03",  x"01",  x"00", -- 0300
         x"00",  x"00",  x"00",  x"00",  x"00",  x"71",  x"fd",  x"77", -- 0308
         x"6e",  x"36",  x"1b",  x"0d",  x"06",  x"80",  x"00",  x"00", -- 0310
         x"00",  x"00",  x"00",  x"80",  x"f0",  x"00",  x"03",  x"07", -- 0318
         x"03",  x"04",  x"04",  x"04",  x"02",  x"c0",  x"e0",  x"c0", -- 0320
         x"40",  x"40",  x"20",  x"20",  x"10",  x"02",  x"02",  x"01", -- 0328
         x"01",  x"01",  x"01",  x"01",  x"01",  x"00",  x"00",  x"00", -- 0330
         x"00",  x"00",  x"00",  x"e0",  x"cc",  x"ff",  x"7f",  x"3d", -- 0338
         x"1e",  x"1e",  x"0f",  x"0e",  x"1c",  x"80",  x"c0",  x"e0", -- 0340
         x"f0",  x"78",  x"78",  x"70",  x"e0",  x"10",  x"08",  x"08", -- 0348
         x"04",  x"04",  x"02",  x"0f",  x"02",  x"33",  x"0c",  x"03", -- 0350
         x"00",  x"00",  x"00",  x"00",  x"00",  x"70",  x"f9",  x"37", -- 0358
         x"ff",  x"3b",  x"0c",  x"03",  x"00",  x"c0",  x"80",  x"00", -- 0360
         x"00",  x"80",  x"c0",  x"33",  x"cc",  x"00",  x"00",  x"1f", -- 0368
         x"3f",  x"7f",  x"ff",  x"00",  x"ff",  x"00",  x"00",  x"ff", -- 0370
         x"7f",  x"7f",  x"7f",  x"ff",  x"ff",  x"00",  x"00",  x"ff", -- 0378
         x"fe",  x"fe",  x"fe",  x"fe",  x"ff",  x"00",  x"00",  x"f8", -- 0380
         x"fc",  x"fe",  x"ff",  x"00",  x"ff",  x"ff",  x"ff",  x"fc", -- 0388
         x"f8",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"3f", -- 0390
         x"1f",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"fc", -- 0398
         x"f8",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"3f", -- 03A0
         x"1f",  x"00",  x"00",  x"00",  x"00",  x"19",  x"ff",  x"ff", -- 03A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
