library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom2_3400 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom2_3400;

architecture rtl of rom2_3400 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"20",  x"45",  x"52",  x"20",  x"57",  x"49",  x"4c",  x"4c", -- 0000
         x"20",  x"49",  x"48",  x"4e",  x"20",  x"20",  x"20",  x"20", -- 0008
         x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20", -- 0010
         x"41",  x"55",  x"46",  x"46",  x"52",  x"45",  x"53",  x"53", -- 0018
         x"45",  x"4e",  x"20",  x"21",  x"20",  x"20",  x"5a",  x"45", -- 0020
         x"49",  x"54",  x"20",  x"3d",  x"20",  x"30",  x"30",  x"3a", -- 0028
         x"20",  x"2d",  x"20",  x"31",  x"20",  x"48",  x"41",  x"53", -- 0030
         x"45",  x"00",  x"50",  x"55",  x"4e",  x"4b",  x"54",  x"45", -- 0038
         x"42",  x"45",  x"57",  x"45",  x"52",  x"54",  x"55",  x"4e", -- 0040
         x"47",  x"3a",  x"20",  x"45",  x"52",  x"42",  x"53",  x"45", -- 0048
         x"3a",  x"20",  x"31",  x"20",  x"50",  x"55",  x"4e",  x"4b", -- 0050
         x"54",  x"20",  x"20",  x"4d",  x"4f",  x"45",  x"48",  x"52", -- 0058
         x"45",  x"3a",  x"20",  x"35",  x"20",  x"50",  x"55",  x"4e", -- 0060
         x"4b",  x"54",  x"45",  x"20",  x"42",  x"49",  x"52",  x"4e", -- 0068
         x"45",  x"3a",  x"20",  x"37",  x"20",  x"42",  x"5a",  x"57", -- 0070
         x"2e",  x"20",  x"31",  x"30",  x"20",  x"50",  x"55",  x"4e", -- 0078
         x"4b",  x"54",  x"45",  x"20",  x"20",  x"2a",  x"20",  x"45", -- 0080
         x"4e",  x"44",  x"45",  x"20",  x"44",  x"45",  x"53",  x"20", -- 0088
         x"53",  x"50",  x"49",  x"45",  x"4c",  x"45",  x"53",  x"20", -- 0090
         x"2a",  x"20",  x"3d",  x"3d",  x"20",  x"52",  x"45",  x"43", -- 0098
         x"4f",  x"52",  x"44",  x"3a",  x"3d",  x"3d",  x"3d",  x"3d", -- 00A0
         x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"20",  x"50",  x"55", -- 00A8
         x"4e",  x"4b",  x"54",  x"45",  x"3a",  x"3d",  x"3d",  x"3d", -- 00B0
         x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"20",  x"48", -- 00B8
         x"41",  x"53",  x"45",  x"4e",  x"3a",  x"3d",  x"3d",  x"3d", -- 00C0
         x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"20", -- 00C8
         x"5a",  x"45",  x"49",  x"54",  x"3a",  x"3d",  x"3d",  x"3d", -- 00D0
         x"3d",  x"3d",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 00D8
         x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 00E0
         x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 00E8
         x"df",  x"df",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00F0
         x"00",  x"00",  x"00",  x"df",  x"df",  x"df",  x"df",  x"df", -- 00F8
         x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 0100
         x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 0108
         x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 0110
         x"df",  x"df",  x"df",  x"e8",  x"e1",  x"00",  x"e8",  x"e1", -- 0118
         x"00",  x"e8",  x"e1",  x"00",  x"e8",  x"e1",  x"00",  x"e8", -- 0120
         x"e1",  x"00",  x"e3",  x"e2",  x"00",  x"e8",  x"e1",  x"00", -- 0128
         x"e8",  x"e1",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0130
         x"00",  x"00",  x"00",  x"df",  x"e8",  x"e1",  x"00",  x"e8", -- 0138
         x"e1",  x"00",  x"e8",  x"e1",  x"00",  x"e8",  x"e1",  x"00", -- 0140
         x"e8",  x"e1",  x"00",  x"e8",  x"e1",  x"00",  x"e3",  x"e2", -- 0148
         x"00",  x"e8",  x"e1",  x"00",  x"e8",  x"e1",  x"00",  x"e8", -- 0150
         x"e1",  x"df",  x"df",  x"e0",  x"e9",  x"00",  x"e0",  x"e9", -- 0158
         x"00",  x"e0",  x"e9",  x"00",  x"e0",  x"e9",  x"00",  x"e0", -- 0160
         x"e9",  x"00",  x"e5",  x"e4",  x"00",  x"e0",  x"e9",  x"00", -- 0168
         x"e0",  x"e9",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0170
         x"00",  x"00",  x"00",  x"df",  x"e0",  x"e9",  x"00",  x"e0", -- 0178
         x"e9",  x"00",  x"e0",  x"e9",  x"00",  x"e0",  x"e9",  x"00", -- 0180
         x"e0",  x"e9",  x"00",  x"e0",  x"e9",  x"00",  x"e5",  x"e4", -- 0188
         x"00",  x"e0",  x"e9",  x"00",  x"e0",  x"e9",  x"00",  x"e0", -- 0190
         x"e9",  x"df",  x"df",  x"00",  x"00",  x"df",  x"df",  x"df", -- 0198
         x"df",  x"df",  x"df",  x"df",  x"00",  x"00",  x"df",  x"df", -- 01A0
         x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 01A8
         x"00",  x"00",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 01B0
         x"df",  x"df",  x"df",  x"df",  x"00",  x"00",  x"df",  x"df", -- 01B8
         x"df",  x"df",  x"df",  x"df",  x"df",  x"00",  x"00",  x"df", -- 01C0
         x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 01C8
         x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"00", -- 01D0
         x"00",  x"df",  x"df",  x"e8",  x"e1",  x"df",  x"00",  x"00", -- 01D8
         x"00",  x"00",  x"00",  x"df",  x"e8",  x"e1",  x"00",  x"e8", -- 01E0
         x"e1",  x"00",  x"e8",  x"e1",  x"00",  x"e8",  x"e1",  x"00", -- 01E8
         x"e8",  x"e1",  x"00",  x"e8",  x"e1",  x"00",  x"e8",  x"e1", -- 01F0
         x"00",  x"e8",  x"e1",  x"00",  x"e8",  x"e1",  x"df",  x"00", -- 01F8
         x"00",  x"00",  x"00",  x"00",  x"df",  x"e8",  x"e1",  x"df", -- 0200
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0208
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"e8", -- 0210
         x"e1",  x"df",  x"df",  x"e0",  x"e9",  x"df",  x"00",  x"00", -- 0218
         x"00",  x"00",  x"00",  x"df",  x"e0",  x"e9",  x"00",  x"e0", -- 0220
         x"e9",  x"00",  x"e0",  x"e9",  x"00",  x"e0",  x"e9",  x"00", -- 0228
         x"e0",  x"e9",  x"00",  x"e0",  x"e9",  x"00",  x"e0",  x"e9", -- 0230
         x"00",  x"e0",  x"e9",  x"00",  x"e0",  x"e9",  x"df",  x"00", -- 0238
         x"00",  x"00",  x"00",  x"00",  x"df",  x"e0",  x"e9",  x"df", -- 0240
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0248
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"e0", -- 0250
         x"e9",  x"df",  x"df",  x"00",  x"00",  x"df",  x"00",  x"00", -- 0258
         x"00",  x"00",  x"00",  x"df",  x"00",  x"00",  x"df",  x"df", -- 0260
         x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 0268
         x"00",  x"00",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 0270
         x"df",  x"df",  x"df",  x"df",  x"00",  x"00",  x"df",  x"00", -- 0278
         x"00",  x"00",  x"00",  x"00",  x"df",  x"00",  x"00",  x"df", -- 0280
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0288
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 0290
         x"00",  x"df",  x"df",  x"e8",  x"e1",  x"df",  x"00",  x"00", -- 0298
         x"00",  x"00",  x"00",  x"df",  x"e8",  x"e1",  x"df",  x"00", -- 02A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df", -- 02A8
         x"e8",  x"e1",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02B0
         x"00",  x"00",  x"00",  x"df",  x"e8",  x"e1",  x"df",  x"00", -- 02B8
         x"00",  x"00",  x"00",  x"00",  x"df",  x"e8",  x"e1",  x"df", -- 02C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"e8", -- 02D0
         x"e1",  x"df",  x"df",  x"e0",  x"e9",  x"df",  x"00",  x"00", -- 02D8
         x"00",  x"00",  x"00",  x"df",  x"e0",  x"e9",  x"df",  x"00", -- 02E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df", -- 02E8
         x"e0",  x"e9",  x"df",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02F0
         x"00",  x"00",  x"00",  x"df",  x"e0",  x"e9",  x"df",  x"00", -- 02F8
         x"00",  x"00",  x"00",  x"00",  x"df",  x"e0",  x"e9",  x"df", -- 0300
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0308
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"e0", -- 0310
         x"e9",  x"df",  x"df",  x"00",  x"00",  x"df",  x"df",  x"df", -- 0318
         x"df",  x"df",  x"df",  x"df",  x"00",  x"00",  x"df",  x"00", -- 0320
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df", -- 0328
         x"00",  x"00",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 0330
         x"df",  x"df",  x"df",  x"df",  x"00",  x"00",  x"df",  x"00", -- 0338
         x"00",  x"00",  x"00",  x"00",  x"df",  x"00",  x"00",  x"df", -- 0340
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0348
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"00", -- 0350
         x"00",  x"00",  x"00",  x"e8",  x"e1",  x"00",  x"e8",  x"e1", -- 0358
         x"00",  x"e8",  x"e1",  x"00",  x"e8",  x"e1",  x"df",  x"00", -- 0360
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df", -- 0368
         x"e8",  x"e1",  x"de",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0370
         x"00",  x"00",  x"00",  x"df",  x"e8",  x"e1",  x"df",  x"00", -- 0378
         x"00",  x"00",  x"00",  x"00",  x"df",  x"e8",  x"e1",  x"df", -- 0380
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0388
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"e8", -- 0390
         x"e1",  x"00",  x"00",  x"e0",  x"e9",  x"00",  x"e0",  x"e9", -- 0398
         x"00",  x"e0",  x"e9",  x"00",  x"e0",  x"e9",  x"df",  x"00", -- 03A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df", -- 03A8
         x"e0",  x"e9",  x"de",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03B0
         x"00",  x"00",  x"00",  x"df",  x"e0",  x"e9",  x"df",  x"00", -- 03B8
         x"00",  x"00",  x"00",  x"00",  x"df",  x"e0",  x"e9",  x"df", -- 03C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"df",  x"e0", -- 03D0
         x"e9",  x"df",  x"df",  x"00",  x"00",  x"df",  x"df",  x"df", -- 03D8
         x"df",  x"df",  x"df",  x"df",  x"00",  x"00",  x"df",  x"df", -- 03E0
         x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 03E8
         x"00",  x"00",  x"df",  x"df",  x"df",  x"df",  x"df",  x"df", -- 03F0
         x"df",  x"df",  x"df",  x"df",  x"00",  x"00",  x"df",  x"df"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
