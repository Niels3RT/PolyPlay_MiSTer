library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_6400 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_6400;

architecture rtl of rom1_6400 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"0d",  x"b7",  x"28",  x"50",  x"ed",  x"52",  x"e5",  x"21", -- 0000
         x"00",  x"0d",  x"36",  x"00",  x"dd",  x"7e",  x"02",  x"c6", -- 0008
         x"04",  x"e6",  x"0e",  x"dd",  x"77",  x"02",  x"cd",  x"c8", -- 0010
         x"66",  x"cd",  x"de",  x"66",  x"e1",  x"19",  x"cd",  x"3f", -- 0018
         x"66",  x"3a",  x"00",  x"0d",  x"b7",  x"28",  x"2d",  x"ed", -- 0020
         x"52",  x"e5",  x"dd",  x"7e",  x"02",  x"3d",  x"3d",  x"e6", -- 0028
         x"0e",  x"dd",  x"77",  x"02",  x"cd",  x"c8",  x"66",  x"cd", -- 0030
         x"e3",  x"66",  x"e1",  x"3a",  x"16",  x"0d",  x"b7",  x"20", -- 0038
         x"19",  x"cd",  x"7f",  x"65",  x"e5",  x"21",  x"d4",  x"68", -- 0040
         x"cd",  x"d4",  x"01",  x"dd",  x"36",  x"03",  x"40",  x"dd", -- 0048
         x"36",  x"04",  x"ff",  x"e1",  x"cd",  x"7f",  x"65",  x"c3", -- 0050
         x"03",  x"62",  x"3e",  x"38",  x"dd",  x"ae",  x"01",  x"dd", -- 0058
         x"77",  x"01",  x"18",  x"f0",  x"ed",  x"52",  x"e5",  x"dd", -- 0060
         x"7e",  x"02",  x"18",  x"c8",  x"3a",  x"bf",  x"0c",  x"47", -- 0068
         x"3e",  x"50",  x"90",  x"4f",  x"32",  x"3d",  x"0c",  x"21", -- 0070
         x"30",  x"f8",  x"22",  x"3f",  x"0c",  x"cd",  x"70",  x"02", -- 0078
         x"36",  x"45",  x"2b",  x"36",  x"53",  x"3a",  x"13",  x"0d", -- 0080
         x"47",  x"cb",  x"21",  x"21",  x"90",  x"65",  x"af",  x"ed", -- 0088
         x"42",  x"4f",  x"57",  x"5f",  x"44",  x"eb",  x"19",  x"30", -- 0090
         x"01",  x"0c",  x"10",  x"fa",  x"41",  x"4c",  x"21",  x"2d", -- 0098
         x"0d",  x"cb",  x"46",  x"28",  x"04",  x"cb",  x"38",  x"cb", -- 00A0
         x"19",  x"21",  x"16",  x"0d",  x"cb",  x"46",  x"28",  x"04", -- 00A8
         x"cb",  x"38",  x"cb",  x"19",  x"cb",  x"38",  x"cb",  x"19", -- 00B0
         x"21",  x"1e",  x"f8",  x"22",  x"3f",  x"0c",  x"2a",  x"18", -- 00B8
         x"0c",  x"09",  x"22",  x"3d",  x"0c",  x"22",  x"18",  x"0c", -- 00C0
         x"cd",  x"70",  x"02",  x"21",  x"c0",  x"f8",  x"3e",  x"0d", -- 00C8
         x"cd",  x"bc",  x"01",  x"cd",  x"72",  x"66",  x"70",  x"67", -- 00D0
         x"21",  x"2d",  x"0d",  x"cb",  x"4e",  x"20",  x"05",  x"21", -- 00D8
         x"21",  x"f9",  x"36",  x"32",  x"cd",  x"72",  x"66",  x"84", -- 00E0
         x"67",  x"21",  x"94",  x"f9",  x"dd",  x"36",  x"00",  x"8e", -- 00E8
         x"cd",  x"7f",  x"65",  x"cd",  x"72",  x"66",  x"8f",  x"67", -- 00F0
         x"21",  x"16",  x"0d",  x"3e",  x"01",  x"ae",  x"77",  x"21", -- 00F8
         x"d4",  x"fa",  x"cd",  x"7f",  x"65",  x"e1",  x"21",  x"2d", -- 0100
         x"0d",  x"3a",  x"16",  x"0d",  x"b7",  x"28",  x"0a",  x"cb", -- 0108
         x"86",  x"21",  x"da",  x"68",  x"cd",  x"e0",  x"01",  x"18", -- 0110
         x"06",  x"21",  x"eb",  x"68",  x"cd",  x"e0",  x"01",  x"06", -- 0118
         x"03",  x"cd",  x"f8",  x"66",  x"21",  x"2d",  x"0d",  x"cb", -- 0120
         x"4e",  x"28",  x"05",  x"cb",  x"8e",  x"c3",  x"34",  x"60", -- 0128
         x"af",  x"32",  x"03",  x"0c",  x"2a",  x"10",  x"0c",  x"ed", -- 0130
         x"4b",  x"18",  x"0c",  x"b7",  x"ed",  x"42",  x"30",  x"04", -- 0138
         x"ed",  x"43",  x"10",  x"0c",  x"fd",  x"77",  x"00",  x"c3", -- 0140
         x"f1",  x"00",  x"21",  x"80",  x"fb",  x"01",  x"40",  x"01", -- 0148
         x"36",  x"8b",  x"23",  x"0b",  x"78",  x"b1",  x"20",  x"f8", -- 0150
         x"cd",  x"72",  x"66",  x"9a",  x"67",  x"21",  x"c3",  x"68", -- 0158
         x"cd",  x"e0",  x"01",  x"18",  x"ba",  x"47",  x"3a",  x"16", -- 0160
         x"0d",  x"b7",  x"78",  x"28",  x"4d",  x"06",  x"01",  x"cd", -- 0168
         x"bc",  x"65",  x"c6",  x"07",  x"06",  x"02",  x"cd",  x"bc", -- 0170
         x"65",  x"d6",  x"07",  x"06",  x"01",  x"18",  x"3d",  x"e5", -- 0178
         x"d5",  x"c5",  x"3a",  x"16",  x"0d",  x"b7",  x"20",  x"18", -- 0180
         x"e5",  x"3e",  x"fd",  x"11",  x"17",  x"0d",  x"cd",  x"54", -- 0188
         x"66",  x"01",  x"3c",  x"00",  x"09",  x"cd",  x"54",  x"66", -- 0190
         x"01",  x"3c",  x"00",  x"09",  x"cd",  x"54",  x"66",  x"e1", -- 0198
         x"dd",  x"7e",  x"01",  x"dd",  x"86",  x"00",  x"0e",  x"01", -- 01A0
         x"11",  x"3c",  x"00",  x"cd",  x"ba",  x"65",  x"19",  x"cd", -- 01A8
         x"65",  x"65",  x"19",  x"cd",  x"ba",  x"65",  x"c1",  x"d1", -- 01B0
         x"e1",  x"c9",  x"06",  x"04",  x"fe",  x"00",  x"20",  x"1b", -- 01B8
         x"cb",  x"7e",  x"28",  x"17",  x"3a",  x"15",  x"0d",  x"be", -- 01C0
         x"3e",  x"00",  x"38",  x"15",  x"3e",  x"f9",  x"be",  x"3e", -- 01C8
         x"00",  x"38",  x"09",  x"3e",  x"80",  x"32",  x"00",  x"0d", -- 01D0
         x"af",  x"18",  x"01",  x"77",  x"23",  x"81",  x"10",  x"dc", -- 01D8
         x"c9",  x"e5",  x"f5",  x"3a",  x"16",  x"0d",  x"b7",  x"20", -- 01E0
         x"06",  x"21",  x"d7",  x"68",  x"cd",  x"d4",  x"01",  x"f1", -- 01E8
         x"21",  x"00",  x"0d",  x"36",  x"01",  x"e1",  x"18",  x"e4", -- 01F0
         x"e5",  x"d5",  x"c5",  x"0e",  x"00",  x"3e",  x"20",  x"18", -- 01F8
         x"a7",  x"e5",  x"d5",  x"c5",  x"f5",  x"3a",  x"16",  x"0d", -- 0200
         x"b7",  x"20",  x"2f",  x"2a",  x"2f",  x"0d",  x"7d",  x"b4", -- 0208
         x"28",  x"15",  x"0e",  x"fd",  x"dd",  x"e5",  x"dd",  x"2a", -- 0210
         x"31",  x"0d",  x"cd",  x"90",  x"66",  x"dd",  x"e1",  x"20", -- 0218
         x"06",  x"21",  x"00",  x"00",  x"22",  x"2f",  x"0d",  x"21", -- 0220
         x"17",  x"0d",  x"5e",  x"23",  x"56",  x"23",  x"7b",  x"b2", -- 0228
         x"28",  x"05",  x"3e",  x"fd",  x"12",  x"18",  x"f3",  x"cd", -- 0230
         x"49",  x"66",  x"f1",  x"c1",  x"d1",  x"e1",  x"c9",  x"e5", -- 0238
         x"d5",  x"c5",  x"0e",  x"00",  x"3e",  x"00",  x"c3",  x"a8", -- 0240
         x"65",  x"21",  x"17",  x"0d",  x"06",  x"14",  x"36",  x"00", -- 0248
         x"23",  x"10",  x"fb",  x"c9",  x"06",  x"04",  x"be",  x"20", -- 0250
         x"06",  x"eb",  x"73",  x"23",  x"72",  x"23",  x"eb",  x"23", -- 0258
         x"10",  x"f4",  x"c9",  x"f5",  x"dd",  x"7e",  x"03",  x"c6", -- 0260
         x"02",  x"fe",  x"40",  x"30",  x"03",  x"dd",  x"77",  x"03", -- 0268
         x"f1",  x"c9",  x"e1",  x"5e",  x"23",  x"56",  x"23",  x"e5", -- 0270
         x"d5",  x"e1",  x"5e",  x"23",  x"56",  x"23",  x"4e",  x"06", -- 0278
         x"00",  x"23",  x"ed",  x"b0",  x"c9",  x"eb",  x"c5",  x"4e", -- 0280
         x"23",  x"06",  x"00",  x"ed",  x"b0",  x"eb",  x"c1",  x"c9", -- 0288
         x"dd",  x"46",  x"00",  x"dd",  x"23",  x"78",  x"b7",  x"c8", -- 0290
         x"dd",  x"7e",  x"00",  x"e5",  x"21",  x"13",  x"69",  x"85", -- 0298
         x"6f",  x"30",  x"01",  x"24",  x"5e",  x"23",  x"56",  x"e1", -- 02A0
         x"19",  x"cb",  x"7e",  x"20",  x"07",  x"71",  x"10",  x"f8", -- 02A8
         x"dd",  x"23",  x"18",  x"dc",  x"3e",  x"fc",  x"be",  x"38", -- 02B0
         x"f4",  x"79",  x"fe",  x"fd",  x"c0",  x"0e",  x"20",  x"dd", -- 02B8
         x"2a",  x"31",  x"0d",  x"2a",  x"2f",  x"0d",  x"18",  x"c8", -- 02C0
         x"21",  x"13",  x"69",  x"85",  x"6f",  x"30",  x"01",  x"24", -- 02C8
         x"5e",  x"23",  x"56",  x"c9",  x"21",  x"01",  x"fc",  x"06", -- 02D0
         x"09",  x"71",  x"23",  x"10",  x"fc",  x"c9",  x"3a",  x"16", -- 02D8
         x"0d",  x"b7",  x"c8",  x"dd",  x"7e",  x"02",  x"21",  x"03", -- 02E0
         x"69",  x"85",  x"6f",  x"30",  x"01",  x"24",  x"7e",  x"dd", -- 02E8
         x"77",  x"00",  x"23",  x"dd",  x"7e",  x"01",  x"be",  x"c9", -- 02F0
         x"3e",  x"4d",  x"32",  x"bf",  x"0c",  x"3a",  x"bf",  x"0c", -- 02F8
         x"b7",  x"20",  x"fa",  x"10",  x"f3",  x"c9",  x"3a",  x"16", -- 0300
         x"0d",  x"b7",  x"c8",  x"21",  x"d3",  x"69",  x"3a",  x"33", -- 0308
         x"0d",  x"c6",  x"04",  x"fe",  x"19",  x"d0",  x"32",  x"33", -- 0310
         x"0d",  x"85",  x"6f",  x"30",  x"01",  x"24",  x"56",  x"2b", -- 0318
         x"5e",  x"2b",  x"ed",  x"53",  x"31",  x"0d",  x"56",  x"2b", -- 0320
         x"5e",  x"ed",  x"53",  x"2f",  x"0d",  x"c9",  x"00",  x"f8", -- 0328
         x"3f",  x"3d",  x"3d",  x"3d",  x"20",  x"52",  x"45",  x"4b", -- 0330
         x"4f",  x"52",  x"44",  x"3a",  x"20",  x"30",  x"30",  x"20", -- 0338
         x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"20",  x"50", -- 0340
         x"55",  x"4e",  x"4b",  x"54",  x"45",  x"3a",  x"20",  x"30", -- 0348
         x"30",  x"20",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"20", -- 0350
         x"5a",  x"45",  x"49",  x"54",  x"3a",  x"20",  x"30",  x"30", -- 0358
         x"2c",  x"30",  x"30",  x"20",  x"53",  x"45",  x"4b",  x"2e", -- 0360
         x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d", -- 0368
         x"18",  x"f9",  x"11",  x"45",  x"52",  x"47",  x"45",  x"42", -- 0370
         x"4e",  x"49",  x"53",  x"20",  x"31",  x"2e",  x"52",  x"45", -- 0378
         x"4e",  x"4e",  x"45",  x"4e",  x"c8",  x"f9",  x"08",  x"31", -- 0380
         x"2e",  x"50",  x"4c",  x"41",  x"54",  x"5a",  x"3a",  x"08", -- 0388
         x"fb",  x"08",  x"32",  x"2e",  x"50",  x"4c",  x"41",  x"54", -- 0390
         x"5a",  x"3a",  x"10",  x"fc",  x"1a",  x"5a",  x"45",  x"49", -- 0398
         x"54",  x"4c",  x"49",  x"4d",  x"49",  x"54",  x"20",  x"55", -- 03A0
         x"45",  x"42",  x"45",  x"52",  x"53",  x"43",  x"48",  x"52", -- 03A8
         x"49",  x"54",  x"54",  x"45",  x"4e",  x"20",  x"21",  x"d2", -- 03B0
         x"f8",  x"08",  x"31",  x"2e",  x"52",  x"45",  x"4e",  x"4e", -- 03B8
         x"45",  x"4e",  x"52",  x"f9",  x"07",  x"31",  x"2e",  x"52", -- 03C0
         x"55",  x"4e",  x"44",  x"45",  x"12",  x"f9",  x"19",  x"4b", -- 03C8
         x"20",  x"2d",  x"20",  x"57",  x"20",  x"41",  x"20",  x"47", -- 03D0
         x"20",  x"45",  x"20",  x"4e",  x"20",  x"52",  x"20",  x"45", -- 03D8
         x"20",  x"4e",  x"20",  x"4e",  x"20",  x"45",  x"20",  x"4e", -- 03E0
         x"89",  x"fa",  x"31",  x"2d",  x"20",  x"48",  x"41",  x"4e", -- 03E8
         x"44",  x"47",  x"45",  x"53",  x"54",  x"45",  x"55",  x"45", -- 03F0
         x"52",  x"54",  x"20",  x"28",  x"47",  x"45",  x"53",  x"43"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
