library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_7800 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_7800;

architecture rtl of rom1_7800 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"c5",  x"47",  x"3e",  x"5d",  x"90",  x"c1",  x"05",  x"28", -- 0000
         x"0f",  x"cb",  x"41",  x"28",  x"1e",  x"19",  x"36",  x"fb", -- 0008
         x"23",  x"36",  x"fb",  x"3d",  x"28",  x"2b",  x"10",  x"f5", -- 0010
         x"dd",  x"23",  x"dd",  x"23",  x"dd",  x"23",  x"dd",  x"46", -- 0018
         x"00",  x"dd",  x"5e",  x"01",  x"dd",  x"56",  x"02",  x"cb", -- 0020
         x"38",  x"30",  x"e2",  x"19",  x"36",  x"fa",  x"11",  x"40", -- 0028
         x"00",  x"19",  x"36",  x"fa",  x"dd",  x"5e",  x"01",  x"dd", -- 0030
         x"56",  x"02",  x"3d",  x"28",  x"04",  x"10",  x"ec",  x"18", -- 0038
         x"d7",  x"c1",  x"d1",  x"e1",  x"dd",  x"e1",  x"c9",  x"dd", -- 0040
         x"21",  x"63",  x"7a",  x"21",  x"ff",  x"7c",  x"47",  x"04", -- 0048
         x"dd",  x"23",  x"dd",  x"23",  x"23",  x"23",  x"23",  x"10", -- 0050
         x"f7",  x"c9",  x"c5",  x"e5",  x"ed",  x"5f",  x"e6",  x"0f", -- 0058
         x"fe",  x"0c",  x"38",  x"03",  x"07",  x"e6",  x"07",  x"e6", -- 0060
         x"0e",  x"47",  x"0f",  x"80",  x"5f",  x"16",  x"00",  x"21", -- 0068
         x"02",  x"7d",  x"19",  x"eb",  x"e1",  x"78",  x"07",  x"c6", -- 0070
         x"80",  x"c1",  x"c9",  x"e5",  x"d5",  x"c5",  x"21",  x"2d", -- 0078
         x"0d",  x"3a",  x"bf",  x"0c",  x"e6",  x"08",  x"be",  x"c4", -- 0080
         x"69",  x"79",  x"3a",  x"bf",  x"0c",  x"b7",  x"c2",  x"18", -- 0088
         x"79",  x"3e",  x"4d",  x"32",  x"bf",  x"0c",  x"21",  x"00", -- 0090
         x"0d",  x"35",  x"7e",  x"32",  x"3d",  x"0c",  x"21",  x"32", -- 0098
         x"f8",  x"22",  x"3f",  x"0c",  x"cd",  x"70",  x"02",  x"2b", -- 00A0
         x"11",  x"f9",  x"7c",  x"cd",  x"68",  x"77",  x"cd",  x"a8", -- 00A8
         x"77",  x"3a",  x"00",  x"0d",  x"fe",  x"06",  x"30",  x"12", -- 00B0
         x"3e",  x"3e",  x"32",  x"60",  x"0c",  x"c6",  x"05",  x"32", -- 00B8
         x"61",  x"0c",  x"3e",  x"55",  x"32",  x"5a",  x"0c",  x"3a", -- 00C0
         x"00",  x"0d",  x"b7",  x"20",  x"4c",  x"21",  x"80",  x"fa", -- 00C8
         x"36",  x"ff",  x"11",  x"81",  x"fa",  x"01",  x"bf",  x"02", -- 00D0
         x"ed",  x"b0",  x"06",  x"05",  x"21",  x"48",  x"fb",  x"11", -- 00D8
         x"10",  x"00",  x"c5",  x"06",  x"30",  x"36",  x"20",  x"23", -- 00E0
         x"10",  x"fb",  x"19",  x"c1",  x"10",  x"f4",  x"cd",  x"55", -- 00E8
         x"77",  x"38",  x"7b",  x"21",  x"38",  x"7d",  x"cd",  x"e0", -- 00F0
         x"01",  x"ed",  x"7b",  x"2b",  x"0d",  x"af",  x"32",  x"03", -- 00F8
         x"0c",  x"fd",  x"77",  x"00",  x"2a",  x"12",  x"0c",  x"ed", -- 0100
         x"4b",  x"18",  x"0c",  x"b7",  x"ed",  x"42",  x"d2",  x"f1", -- 0108
         x"00",  x"ed",  x"43",  x"12",  x"0c",  x"c3",  x"f1",  x"00", -- 0110
         x"af",  x"c1",  x"d1",  x"e1",  x"c9",  x"e5",  x"2a",  x"27", -- 0118
         x"0d",  x"22",  x"3d",  x"0c",  x"21",  x"f0",  x"fc",  x"22", -- 0120
         x"3f",  x"0c",  x"cd",  x"70",  x"02",  x"36",  x"20",  x"2b", -- 0128
         x"36",  x"20",  x"af",  x"2a",  x"27",  x"0d",  x"11",  x"1e", -- 0130
         x"00",  x"3c",  x"ed",  x"52",  x"30",  x"fb",  x"fe",  x"3d", -- 0138
         x"38",  x"02",  x"3e",  x"3c",  x"32",  x"29",  x"0d",  x"32", -- 0140
         x"3d",  x"0c",  x"21",  x"f0",  x"fd",  x"22",  x"3f",  x"0c", -- 0148
         x"cd",  x"70",  x"02",  x"36",  x"20",  x"2b",  x"36",  x"20", -- 0150
         x"e1",  x"c9",  x"f5",  x"cd",  x"d4",  x"01",  x"cd",  x"7b", -- 0158
         x"78",  x"3a",  x"59",  x"0c",  x"b7",  x"20",  x"f7",  x"f1", -- 0160
         x"c9",  x"32",  x"2d",  x"0d",  x"3a",  x"2e",  x"0d",  x"b7", -- 0168
         x"c8",  x"dd",  x"e5",  x"2a",  x"2f",  x"0d",  x"11",  x"18", -- 0170
         x"00",  x"19",  x"e5",  x"dd",  x"e1",  x"3a",  x"2d",  x"0d", -- 0178
         x"b7",  x"28",  x"07",  x"3e",  x"9c",  x"cd",  x"88",  x"77", -- 0180
         x"18",  x"03",  x"cd",  x"81",  x"77",  x"dd",  x"e1",  x"c9", -- 0188
         x"d5",  x"16",  x"20",  x"18",  x"03",  x"d5",  x"16",  x"f8", -- 0190
         x"c5",  x"f5",  x"e5",  x"dd",  x"6e",  x"00",  x"dd",  x"66", -- 0198
         x"01",  x"01",  x"be",  x"ff",  x"09",  x"06",  x"04",  x"23", -- 01A0
         x"72",  x"10",  x"fc",  x"01",  x"40",  x"00",  x"09",  x"72", -- 01A8
         x"09",  x"72",  x"09",  x"06",  x"04",  x"72",  x"2b",  x"10", -- 01B0
         x"fc",  x"23",  x"01",  x"c0",  x"ff",  x"09",  x"72",  x"09", -- 01B8
         x"72",  x"e1",  x"f1",  x"c1",  x"d1",  x"c9",  x"d6",  x"80", -- 01C0
         x"0f",  x"47",  x"0f",  x"80",  x"21",  x"02",  x"7d",  x"85", -- 01C8
         x"6f",  x"30",  x"01",  x"24",  x"cd",  x"95",  x"79",  x"cd", -- 01D0
         x"5a",  x"79",  x"cd",  x"90",  x"79",  x"dd",  x"23",  x"dd", -- 01D8
         x"23",  x"c9",  x"cd",  x"47",  x"78",  x"3e",  x"98",  x"cd", -- 01E0
         x"88",  x"77",  x"3e",  x"80",  x"dd",  x"21",  x"71",  x"7a", -- 01E8
         x"06",  x"06",  x"cd",  x"88",  x"77",  x"3c",  x"10",  x"fa", -- 01F0
         x"c9",  x"cd",  x"7b",  x"78",  x"c8",  x"3a",  x"00",  x"0d", -- 01F8
         x"fe",  x"07",  x"38",  x"0b",  x"e6",  x"07",  x"fe",  x"01", -- 0200
         x"28",  x"0b",  x"fe",  x"04",  x"28",  x"2e",  x"c9",  x"3e", -- 0208
         x"5a",  x"32",  x"00",  x"0d",  x"c9",  x"e5",  x"3e",  x"03", -- 0210
         x"21",  x"00",  x"f9",  x"cd",  x"56",  x"7a",  x"ed",  x"5f", -- 0218
         x"e6",  x"07",  x"c6",  x"03",  x"32",  x"24",  x"0d",  x"47", -- 0220
         x"dd",  x"21",  x"95",  x"7a",  x"cd",  x"5a",  x"78",  x"cd", -- 0228
         x"88",  x"77",  x"21",  x"ff",  x"7c",  x"cd",  x"5a",  x"79", -- 0230
         x"10",  x"f2",  x"e1",  x"c9",  x"e5",  x"3e",  x"03",  x"21", -- 0238
         x"00",  x"f9",  x"cd",  x"56",  x"7a",  x"3a",  x"24",  x"0d", -- 0240
         x"47",  x"dd",  x"21",  x"95",  x"7a",  x"3e",  x"9c",  x"cd", -- 0248
         x"88",  x"77",  x"10",  x"f9",  x"e1",  x"c9",  x"c5",  x"06", -- 0250
         x"3e",  x"23",  x"36",  x"20",  x"23",  x"10",  x"fb",  x"23", -- 0258
         x"3d",  x"c1",  x"20",  x"f2",  x"c9",  x"4b",  x"fb",  x"0b", -- 0260
         x"fc",  x"cb",  x"fc",  x"8b",  x"fd",  x"4b",  x"fe",  x"0b", -- 0268
         x"ff",  x"47",  x"fb",  x"07",  x"fc",  x"c7",  x"fc",  x"87", -- 0270
         x"fd",  x"47",  x"fe",  x"07",  x"ff",  x"cc",  x"f9",  x"d0", -- 0278
         x"f9",  x"d4",  x"f9",  x"d8",  x"f9",  x"dc",  x"f9",  x"e0", -- 0280
         x"f9",  x"e4",  x"f9",  x"e8",  x"f9",  x"ec",  x"f9",  x"f0", -- 0288
         x"f9",  x"f4",  x"f9",  x"f8",  x"f9",  x"0c",  x"f9",  x"10", -- 0290
         x"f9",  x"14",  x"f9",  x"18",  x"f9",  x"1c",  x"f9",  x"20", -- 0298
         x"f9",  x"24",  x"f9",  x"28",  x"f9",  x"2c",  x"f9",  x"30", -- 02A0
         x"f9",  x"34",  x"f9",  x"38",  x"f9",  x"1c",  x"fd",  x"ff", -- 02A8
         x"03",  x"fe",  x"ff",  x"1d",  x"40",  x"00",  x"02",  x"40", -- 02B0
         x"00",  x"3e",  x"01",  x"00",  x"03",  x"80",  x"ff",  x"1d", -- 02B8
         x"40",  x"ff",  x"02",  x"be",  x"ff",  x"20",  x"fd",  x"ff", -- 02C0
         x"1c",  x"fa",  x"00",  x"f8",  x"3f",  x"3d",  x"3d",  x"3d", -- 02C8
         x"20",  x"52",  x"45",  x"4b",  x"4f",  x"52",  x"44",  x"3a", -- 02D0
         x"20",  x"30",  x"30",  x"20",  x"3d",  x"3d",  x"3d",  x"3d", -- 02D8
         x"3d",  x"3d",  x"20",  x"50",  x"55",  x"4e",  x"4b",  x"54", -- 02E0
         x"45",  x"3a",  x"20",  x"30",  x"30",  x"20",  x"3d",  x"3d", -- 02E8
         x"3d",  x"3d",  x"3d",  x"20",  x"53",  x"50",  x"49",  x"45", -- 02F0
         x"4c",  x"5a",  x"45",  x"49",  x"54",  x"3a",  x"20",  x"39", -- 02F8
         x"30",  x"20",  x"53",  x"45",  x"4b",  x"2e",  x"3d",  x"3d", -- 0300
         x"3d",  x"3d",  x"3d",  x"3d",  x"e5",  x"fb",  x"0c",  x"47", -- 0308
         x"45",  x"57",  x"49",  x"4e",  x"4e",  x"43",  x"48",  x"41", -- 0310
         x"4e",  x"43",  x"45",  x"e0",  x"fc",  x"0c",  x"50",  x"55", -- 0318
         x"4e",  x"4b",  x"54",  x"47",  x"45",  x"57",  x"49",  x"4e", -- 0320
         x"4e",  x"3a",  x"e0",  x"fd",  x"0b",  x"5a",  x"45",  x"49", -- 0328
         x"54",  x"47",  x"45",  x"57",  x"49",  x"4e",  x"4e",  x"3a", -- 0330
         x"d1",  x"fb",  x"1e",  x"2a",  x"2a",  x"2a",  x"2a",  x"2a", -- 0338
         x"20",  x"20",  x"45",  x"4e",  x"44",  x"45",  x"20",  x"44", -- 0340
         x"45",  x"53",  x"20",  x"53",  x"50",  x"49",  x"45",  x"4c", -- 0348
         x"45",  x"53",  x"20",  x"20",  x"2a",  x"2a",  x"2a",  x"2a", -- 0350
         x"2a",  x"43",  x"fa",  x"39",  x"2a",  x"2a",  x"2a",  x"20", -- 0358
         x"4e",  x"41",  x"43",  x"48",  x"42",  x"49",  x"4c",  x"44", -- 0360
         x"45",  x"4e",  x"20",  x"44",  x"45",  x"52",  x"20",  x"44", -- 0368
         x"55",  x"52",  x"43",  x"48",  x"20",  x"20",  x"20",  x"20", -- 0370
         x"56",  x"45",  x"52",  x"44",  x"45",  x"43",  x"4b",  x"54", -- 0378
         x"45",  x"4e",  x"20",  x"42",  x"49",  x"4c",  x"44",  x"2d", -- 0380
         x"2f",  x"54",  x"4f",  x"4e",  x"46",  x"4f",  x"4c",  x"47", -- 0388
         x"45",  x"20",  x"2a",  x"2a",  x"2a",  x"50",  x"fb",  x"2f", -- 0390
         x"2d",  x"50",  x"4f",  x"53",  x"49",  x"54",  x"49",  x"4f", -- 0398
         x"4e",  x"49",  x"45",  x"52",  x"45",  x"20",  x"44",  x"45", -- 03A0
         x"4e",  x"20",  x"47",  x"52",  x"55",  x"45",  x"4e",  x"45", -- 03A8
         x"4e",  x"20",  x"50",  x"46",  x"45",  x"49",  x"4c",  x"20", -- 03B0
         x"4d",  x"49",  x"54",  x"20",  x"44",  x"45",  x"4d",  x"20", -- 03B8
         x"53",  x"54",  x"45",  x"55",  x"45",  x"52",  x"2d",  x"91", -- 03C0
         x"fb",  x"21",  x"4b",  x"4e",  x"55",  x"45",  x"50",  x"50", -- 03C8
         x"45",  x"4c",  x"20",  x"28",  x"4e",  x"41",  x"43",  x"48", -- 03D0
         x"20",  x"4f",  x"42",  x"45",  x"4e",  x"20",  x"2f",  x"20", -- 03D8
         x"4e",  x"41",  x"43",  x"48",  x"20",  x"55",  x"4e",  x"54", -- 03E0
         x"45",  x"4e",  x"29",  x"10",  x"fc",  x"28",  x"2d",  x"45", -- 03E8
         x"49",  x"4e",  x"54",  x"52",  x"41",  x"47",  x"45",  x"4e", -- 03F0
         x"20",  x"44",  x"45",  x"53",  x"20",  x"42",  x"49",  x"4c"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
