library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_zre_0000 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_zre_0000;

architecture rtl of rom_zre_0000 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"31",  x"ff",  x"0f",  x"c3",  x"b3",  x"00",  x"48",  x"3a", -- 0000
         x"c9",  x"20",  x"31",  x"20",  x"4c",  x"45",  x"42",  x"45", -- 0008
         x"c9",  x"20",  x"20",  x"3c",  x"3d",  x"3e",  x"20",  x"20", -- 0010
         x"c9",  x"34",  x"20",  x"53",  x"43",  x"48",  x"55",  x"53", -- 0018
         x"c9",  x"00",  x"00",  x"80",  x"20",  x"00",  x"3d",  x"3d", -- 0020
         x"c9",  x"52",  x"45",  x"43",  x"4f",  x"52",  x"44",  x"3a", -- 0028
         x"c9",  x"30",  x"30",  x"30",  x"20",  x"3d",  x"3d",  x"3d", -- 0030
         x"c9",  x"54",  x"52",  x"45",  x"46",  x"46",  x"45",  x"52", -- 0038
         x"3a",  x"30",  x"30",  x"30",  x"30",  x"20",  x"80",  x"20", -- 0040
         x"60",  x"02",  x"60",  x"02",  x"02",  x"08",  x"ea",  x"01", -- 0048
         x"04",  x"08",  x"60",  x"02",  x"4e",  x"3a",  x"30",  x"30", -- 0050
         x"30",  x"20",  x"3d",  x"3d",  x"3d",  x"20",  x"4c",  x"45", -- 0058
         x"42",  x"45",  x"4e",  x"3a",  x"30",  x"30",  x"08",  x"d9", -- 0060
         x"21",  x"62",  x"0c",  x"23",  x"46",  x"23",  x"7e",  x"23", -- 0068
         x"b7",  x"7e",  x"20",  x"06",  x"b7",  x"28",  x"15",  x"35", -- 0070
         x"18",  x"2a",  x"cb",  x"7f",  x"28",  x"04",  x"e6",  x"7f", -- 0078
         x"20",  x"f5",  x"2a",  x"66",  x"0c",  x"7e",  x"3c",  x"20", -- 0080
         x"0f",  x"32",  x"64",  x"0c",  x"21",  x"62",  x"0c",  x"34", -- 0088
         x"7e",  x"e6",  x"03",  x"47",  x"3e",  x"05",  x"18",  x"09", -- 0090
         x"46",  x"23",  x"7e",  x"23",  x"22",  x"66",  x"0c",  x"cb", -- 0098
         x"ff",  x"32",  x"65",  x"0c",  x"78",  x"32",  x"63",  x"0c", -- 00A0
         x"db",  x"85",  x"e6",  x"e8",  x"b0",  x"d3",  x"85",  x"d9", -- 00A8
         x"08",  x"ed",  x"45",  x"21",  x"ff",  x"0f",  x"11",  x"01", -- 00B0
         x"0c",  x"af",  x"ed",  x"52",  x"44",  x"4d",  x"21",  x"00", -- 00B8
         x"0c",  x"77",  x"ed",  x"b0",  x"21",  x"48",  x"00",  x"7d", -- 00C0
         x"d3",  x"80",  x"7c",  x"ed",  x"47",  x"00",  x"00",  x"00", -- 00C8
         x"ed",  x"5e",  x"fb",  x"3e",  x"ff",  x"d3",  x"86",  x"d3", -- 00D0
         x"86",  x"d3",  x"87",  x"3e",  x"18",  x"d3",  x"87",  x"3e", -- 00D8
         x"60",  x"d3",  x"85",  x"21",  x"50",  x"00",  x"7d",  x"d3", -- 00E0
         x"86",  x"3e",  x"a5",  x"d3",  x"83",  x"3e",  x"80",  x"d3", -- 00E8
         x"83",  x"cd",  x"8f",  x"01",  x"cb",  x"77",  x"28",  x"53", -- 00F0
         x"3e",  x"f7",  x"d3",  x"86",  x"3e",  x"7f",  x"d3",  x"86", -- 00F8
         x"cd",  x"00",  x"08",  x"28",  x"0a",  x"21",  x"00",  x"00", -- 0100
         x"22",  x"18",  x"0c",  x"00",  x"00",  x"00",  x"00",  x"78", -- 0108
         x"ee",  x"07",  x"32",  x"02",  x"0c",  x"3c",  x"3d",  x"ca", -- 0110
         x"00",  x"1c",  x"3d",  x"ca",  x"00",  x"28",  x"3d",  x"ca", -- 0118
         x"00",  x"10",  x"3d",  x"ca",  x"00",  x"40",  x"3d",  x"ca", -- 0120
         x"00",  x"50",  x"3d",  x"ca",  x"00",  x"60",  x"3d",  x"ca", -- 0128
         x"00",  x"74",  x"3d",  x"ca",  x"00",  x"80",  x"cd",  x"b7", -- 0130
         x"01",  x"21",  x"e4",  x"02",  x"11",  x"10",  x"fc",  x"01", -- 0138
         x"20",  x"00",  x"ed",  x"b0",  x"cd",  x"9a",  x"01",  x"20", -- 0140
         x"a8",  x"18",  x"f9",  x"cd",  x"b7",  x"01",  x"2a",  x"00", -- 0148
         x"0c",  x"22",  x"3d",  x"0c",  x"21",  x"00",  x"f8",  x"11", -- 0150
         x"dc",  x"03",  x"19",  x"22",  x"3f",  x"0c",  x"cd",  x"70", -- 0158
         x"02",  x"23",  x"23",  x"eb",  x"21",  x"04",  x"03",  x"01", -- 0160
         x"06",  x"00",  x"ed",  x"b0",  x"cd",  x"84",  x"01",  x"cb", -- 0168
         x"77",  x"28",  x"f9",  x"cd",  x"8f",  x"01",  x"cb",  x"77", -- 0170
         x"20",  x"f9",  x"cd",  x"84",  x"01",  x"cb",  x"77",  x"28", -- 0178
         x"f9",  x"c3",  x"f1",  x"00",  x"06",  x"14",  x"0e",  x"ff", -- 0180
         x"db",  x"84",  x"a1",  x"4f",  x"10",  x"fa",  x"c9",  x"06", -- 0188
         x"14",  x"0e",  x"00",  x"db",  x"84",  x"b1",  x"4f",  x"10", -- 0190
         x"fa",  x"c9",  x"cd",  x"8f",  x"01",  x"2f",  x"cb",  x"77", -- 0198
         x"c0",  x"97",  x"c9",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"3e", -- 01B0
         x"20",  x"21",  x"00",  x"f8",  x"06",  x"40",  x"36",  x"00", -- 01B8
         x"23",  x"10",  x"fb",  x"3d",  x"20",  x"f6",  x"c9",  x"3e", -- 01C0
         x"12",  x"4f",  x"3a",  x"56",  x"0c",  x"3d",  x"20",  x"fd", -- 01C8
         x"0d",  x"20",  x"f7",  x"c9",  x"22",  x"5c",  x"0c",  x"3e", -- 01D0
         x"55",  x"32",  x"58",  x"0c",  x"32",  x"59",  x"0c",  x"c9", -- 01D8
         x"cd",  x"d4",  x"01",  x"3a",  x"59",  x"0c",  x"b7",  x"20", -- 01E0
         x"fa",  x"c9",  x"f5",  x"c5",  x"e5",  x"fb",  x"21",  x"bf", -- 01E8
         x"0c",  x"7e",  x"b7",  x"28",  x"01",  x"35",  x"3a",  x"58", -- 01F0
         x"0c",  x"b7",  x"20",  x"10",  x"3a",  x"59",  x"0c",  x"b7", -- 01F8
         x"28",  x"3d",  x"21",  x"5b",  x"0c",  x"7e",  x"b7",  x"28", -- 0200
         x"0d",  x"35",  x"18",  x"33",  x"2a",  x"5c",  x"0c",  x"22", -- 0208
         x"5e",  x"0c",  x"af",  x"32",  x"58",  x"0c",  x"2a",  x"5e", -- 0210
         x"0c",  x"7e",  x"b7",  x"20",  x"0a",  x"af",  x"32",  x"59", -- 0218
         x"0c",  x"3e",  x"41",  x"d3",  x"80",  x"18",  x"18",  x"47", -- 0220
         x"e6",  x"c0",  x"0f",  x"f6",  x"05",  x"d3",  x"80",  x"23", -- 0228
         x"7e",  x"d3",  x"80",  x"78",  x"23",  x"e6",  x"3f",  x"32", -- 0230
         x"5b",  x"0c",  x"22",  x"5e",  x"0c",  x"28",  x"d7",  x"3a", -- 0238
         x"5a",  x"0c",  x"b7",  x"28",  x"18",  x"3e",  x"05",  x"d3", -- 0240
         x"81",  x"3a",  x"60",  x"0c",  x"3c",  x"21",  x"61",  x"0c", -- 0248
         x"be",  x"20",  x"05",  x"af",  x"32",  x"5a",  x"0c",  x"3c", -- 0250
         x"d3",  x"81",  x"32",  x"60",  x"0c",  x"e1",  x"c1",  x"f1", -- 0258
         x"ed",  x"4d",  x"f5",  x"3e",  x"03",  x"d3",  x"86",  x"3e", -- 0260
         x"55",  x"32",  x"03",  x"0c",  x"fb",  x"f1",  x"ed",  x"4d", -- 0268
         x"af",  x"11",  x"10",  x"27",  x"cd",  x"9a",  x"02",  x"11", -- 0270
         x"e8",  x"03",  x"cd",  x"9a",  x"02",  x"11",  x"64",  x"00", -- 0278
         x"cd",  x"9a",  x"02",  x"3e",  x"30",  x"11",  x"0a",  x"00", -- 0280
         x"cd",  x"9a",  x"02",  x"3a",  x"3d",  x"0c",  x"cd",  x"aa", -- 0288
         x"02",  x"36",  x"00",  x"23",  x"36",  x"3d",  x"23",  x"36", -- 0290
         x"3d",  x"c9",  x"b7",  x"2a",  x"3d",  x"0c",  x"ed",  x"52", -- 0298
         x"38",  x"06",  x"22",  x"3d",  x"0c",  x"3c",  x"18",  x"f2", -- 02A0
         x"b7",  x"c8",  x"f6",  x"30",  x"2a",  x"3f",  x"0c",  x"77", -- 02A8
         x"23",  x"22",  x"3f",  x"0c",  x"3e",  x"30",  x"c9",  x"01", -- 02B0
         x"00",  x"14",  x"21",  x"ff",  x"ff",  x"af",  x"77",  x"0b", -- 02B8
         x"2b",  x"b8",  x"20",  x"fa",  x"b9",  x"20",  x"f7",  x"c9", -- 02C0
         x"d5",  x"11",  x"00",  x"f4",  x"18",  x"0c",  x"d5",  x"11", -- 02C8
         x"00",  x"f0",  x"18",  x"06",  x"d5",  x"11",  x"00",  x"ec", -- 02D0
         x"18",  x"00",  x"29",  x"29",  x"29",  x"19",  x"d1",  x"eb", -- 02D8
         x"ed",  x"b0",  x"eb",  x"c9",  x"47",  x"45",  x"57",  x"41", -- 02E0
         x"45",  x"48",  x"4c",  x"54",  x"45",  x"53",  x"20",  x"53", -- 02E8
         x"50",  x"49",  x"45",  x"4c",  x"20",  x"4e",  x"49",  x"43", -- 02F0
         x"48",  x"54",  x"20",  x"56",  x"4f",  x"52",  x"48",  x"41", -- 02F8
         x"4e",  x"44",  x"45",  x"4e",  x"53",  x"50",  x"49",  x"45", -- 0300
         x"4c",  x"45",  x"20",  x"53",  x"50",  x"49",  x"45",  x"4c", -- 0308
         x"42",  x"45",  x"47",  x"49",  x"4e",  x"4e",  x"20",  x"2d", -- 0310
         x"2d",  x"20",  x"47",  x"45",  x"4c",  x"44",  x"45",  x"49", -- 0318
         x"4e",  x"57",  x"55",  x"52",  x"46",  x"20",  x"06",  x"02", -- 0320
         x"0e",  x"ff",  x"18",  x"02",  x"0e",  x"b0",  x"3e",  x"05", -- 0328
         x"d3",  x"80",  x"79",  x"d3",  x"80",  x"cd",  x"6c",  x"03", -- 0330
         x"0d",  x"3e",  x"50",  x"b9",  x"20",  x"f0",  x"21",  x"00", -- 0338
         x"08",  x"2b",  x"7d",  x"b4",  x"20",  x"fb",  x"0e",  x"50", -- 0340
         x"3e",  x"05",  x"d3",  x"80",  x"79",  x"d3",  x"80",  x"cd", -- 0348
         x"6c",  x"03",  x"0c",  x"3e",  x"01",  x"b8",  x"20",  x"04", -- 0350
         x"3e",  x"ff",  x"18",  x"02",  x"3e",  x"b0",  x"b9",  x"20", -- 0358
         x"e7",  x"10",  x"c9",  x"3e",  x"05",  x"d3",  x"80",  x"3e", -- 0360
         x"01",  x"d3",  x"80",  x"c9",  x"1e",  x"05",  x"79",  x"2f", -- 0368
         x"3d",  x"20",  x"fd",  x"1d",  x"20",  x"f8",  x"c9",  x"00", -- 0370
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0378
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0380
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0388
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0390
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0398
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03A0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03A8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03B0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03B8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03C0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03C8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03D0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03D8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03E0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
