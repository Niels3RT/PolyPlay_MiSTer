library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom2_4c00 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom2_4c00;

architecture rtl of rom2_4c00 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"ff",  x"ff",  x"f3",  x"fd",  x"fe",  x"fe",  x"fe",  x"fe", -- 0000
         x"fe",  x"fe",  x"e7",  x"5f",  x"3f",  x"3f",  x"3f",  x"3f", -- 0008
         x"3f",  x"3f",  x"fe",  x"fe",  x"fe",  x"fe",  x"ff",  x"ff", -- 0010
         x"ff",  x"ff",  x"3f",  x"3f",  x"3f",  x"3f",  x"7f",  x"7f", -- 0018
         x"ff",  x"ff",  x"f3",  x"8d",  x"86",  x"92",  x"d8",  x"cc", -- 0020
         x"cc",  x"ec",  x"e7",  x"58",  x"30",  x"24",  x"0d",  x"19", -- 0028
         x"19",  x"1b",  x"ec",  x"ec",  x"d8",  x"80",  x"83",  x"e7", -- 0030
         x"ff",  x"ff",  x"1b",  x"1b",  x"0d",  x"00",  x"60",  x"73", -- 0038
         x"ff",  x"ff",  x"f3",  x"8d",  x"86",  x"92",  x"d8",  x"cc", -- 0040
         x"cc",  x"ec",  x"e7",  x"58",  x"30",  x"24",  x"0d",  x"19", -- 0048
         x"19",  x"1b",  x"ec",  x"ec",  x"d8",  x"80",  x"83",  x"e7", -- 0050
         x"ff",  x"ff",  x"1b",  x"1b",  x"0d",  x"00",  x"60",  x"73", -- 0058
         x"ff",  x"ff",  x"f3",  x"8d",  x"86",  x"82",  x"c0",  x"c0", -- 0060
         x"c0",  x"e0",  x"e7",  x"58",  x"30",  x"20",  x"01",  x"01", -- 0068
         x"01",  x"03",  x"e4",  x"ee",  x"c6",  x"80",  x"83",  x"e7", -- 0070
         x"ff",  x"ff",  x"13",  x"3b",  x"31",  x"00",  x"60",  x"73", -- 0078
         x"ff",  x"ff",  x"f3",  x"dd",  x"a6",  x"d6",  x"c8",  x"e5", -- 0080
         x"c6",  x"f1",  x"e7",  x"5d",  x"32",  x"35",  x"09",  x"4b", -- 0088
         x"19",  x"47",  x"e4",  x"ff",  x"c6",  x"c5",  x"a3",  x"ef", -- 0090
         x"ff",  x"ff",  x"13",  x"7f",  x"31",  x"51",  x"62",  x"7b", -- 0098
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"fe", -- 00A0
         x"ff",  x"4f",  x"ff",  x"f9",  x"f0",  x"e6",  x"d4",  x"18", -- 00A8
         x"00",  x"80",  x"bf",  x"af",  x"3f",  x"1f",  x"0f",  x"07", -- 00B0
         x"0f",  x"0f",  x"07",  x"07",  x"83",  x"c1",  x"f0",  x"f8", -- 00B8
         x"fc",  x"fc",  x"c0",  x"80",  x"80",  x"00",  x"00",  x"00", -- 00C0
         x"00",  x"00",  x"1f",  x"3f",  x"3f",  x"7f",  x"7f",  x"3f", -- 00C8
         x"1f",  x"1f",  x"f8",  x"d0",  x"c0",  x"80",  x"c0",  x"90", -- 00D0
         x"f8",  x"f8",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00D8
         x"00",  x"00",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f", -- 00E0
         x"0f",  x"0f",  x"f8",  x"fc",  x"fe",  x"ff",  x"ff",  x"f0", -- 00E8
         x"e0",  x"ff",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00F0
         x"00",  x"ff",  x"0f",  x"1f",  x"1f",  x"3f",  x"7f",  x"ff", -- 00F8
         x"ff",  x"ff",  x"fd",  x"f5",  x"fc",  x"f8",  x"f0",  x"e0", -- 0100
         x"f0",  x"f0",  x"ff",  x"9f",  x"0f",  x"67",  x"2b",  x"18", -- 0108
         x"00",  x"01",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7f", -- 0110
         x"ff",  x"f2",  x"f8",  x"fc",  x"fc",  x"fe",  x"fe",  x"fc", -- 0118
         x"f8",  x"f8",  x"03",  x"01",  x"01",  x"00",  x"00",  x"00", -- 0120
         x"00",  x"00",  x"e0",  x"e0",  x"c1",  x"83",  x"0f",  x"1f", -- 0128
         x"3f",  x"3f",  x"f0",  x"f0",  x"f0",  x"f0",  x"f0",  x"f0", -- 0130
         x"f0",  x"f0",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0138
         x"00",  x"00",  x"1f",  x"0b",  x"03",  x"01",  x"03",  x"09", -- 0140
         x"1f",  x"1f",  x"f0",  x"f8",  x"f8",  x"fc",  x"fe",  x"ff", -- 0148
         x"ff",  x"ff",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0150
         x"00",  x"ff",  x"1f",  x"3f",  x"7f",  x"ff",  x"ff",  x"0f", -- 0158
         x"07",  x"ff",  x"aa",  x"55",  x"aa",  x"55",  x"aa",  x"55", -- 0160
         x"aa",  x"00",  x"2a",  x"15",  x"2a",  x"15",  x"2a",  x"15", -- 0168
         x"2a",  x"00",  x"0a",  x"05",  x"0a",  x"05",  x"0a",  x"05", -- 0170
         x"0a",  x"00",  x"02",  x"01",  x"02",  x"01",  x"02",  x"01", -- 0178
         x"02",  x"00",  x"fe",  x"f1",  x"ca",  x"39",  x"b9",  x"c6", -- 0180
         x"f7",  x"f9",  x"00",  x"9c",  x"5a",  x"e5",  x"e5",  x"db", -- 0188
         x"3b",  x"37",  x"47",  x"af",  x"df",  x"ef",  x"f7",  x"f9", -- 0190
         x"fe",  x"ff",  x"fc",  x"fa",  x"f5",  x"ed",  x"d3",  x"b8", -- 0198
         x"b7",  x"00",  x"3f",  x"df",  x"6f",  x"a3",  x"9b",  x"1d", -- 01A0
         x"ee",  x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 01A8
         x"ff",  x"00",  x"7f",  x"8f",  x"53",  x"9c",  x"9d",  x"63", -- 01B0
         x"ef",  x"9f",  x"00",  x"39",  x"5a",  x"a7",  x"a7",  x"db", -- 01B8
         x"dc",  x"ec",  x"e2",  x"f5",  x"fb",  x"f7",  x"ef",  x"9f", -- 01C0
         x"7f",  x"ff",  x"3f",  x"5f",  x"af",  x"b7",  x"cb",  x"1d", -- 01C8
         x"ed",  x"00",  x"fc",  x"fb",  x"f6",  x"c5",  x"d9",  x"b8", -- 01D0
         x"77",  x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 01D8
         x"ff",  x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 01E0
         x"ff",  x"ff",  x"f8",  x"02",  x"00",  x"00",  x"00",  x"39", -- 01E8
         x"3d",  x"1f",  x"0f",  x"7f",  x"00",  x"00",  x"80",  x"ce", -- 01F0
         x"de",  x"fc",  x"f8",  x"ff",  x"ff",  x"0f",  x"1f",  x"3d", -- 01F8
         x"39",  x"00",  x"00",  x"00",  x"ff",  x"f8",  x"fc",  x"de", -- 0200
         x"ce",  x"80",  x"00",  x"00",  x"00",  x"00",  x"00",  x"39", -- 0208
         x"3d",  x"1f",  x"0c",  x"78",  x"00",  x"00",  x"80",  x"ce", -- 0210
         x"de",  x"7c",  x"18",  x"0f",  x"f8",  x"0c",  x"1f",  x"3d", -- 0218
         x"39",  x"00",  x"00",  x"00",  x"0f",  x"18",  x"7c",  x"de", -- 0220
         x"ce",  x"80",  x"00",  x"00",  x"00",  x"00",  x"00",  x"39", -- 0228
         x"3d",  x"1f",  x"0f",  x"7f",  x"00",  x"00",  x"80",  x"ce", -- 0230
         x"de",  x"fc",  x"f8",  x"ff",  x"ff",  x"0f",  x"1f",  x"3d", -- 0238
         x"39",  x"00",  x"00",  x"00",  x"ff",  x"f8",  x"fc",  x"de", -- 0240
         x"ce",  x"80",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0248
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0250
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0258
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0260
         x"00",  x"00",  x"00",  x"00",  x"00",  x"70",  x"78",  x"7c", -- 0268
         x"3e",  x"3e",  x"3e",  x"1e",  x"00",  x"07",  x"0f",  x"1f", -- 0270
         x"3e",  x"3e",  x"3e",  x"3c",  x"1e",  x"1e",  x"3e",  x"3e", -- 0278
         x"3c",  x"18",  x"00",  x"00",  x"3c",  x"3c",  x"3e",  x"3f", -- 0280
         x"1f",  x"0c",  x"00",  x"00",  x"a0",  x"00",  x"00",  x"70", -- 0288
         x"78",  x"7c",  x"3e",  x"3e",  x"3e",  x"1e",  x"00",  x"07", -- 0290
         x"0f",  x"1f",  x"3e",  x"3e",  x"3e",  x"3c",  x"1e",  x"1e", -- 0298
         x"3e",  x"3e",  x"3c",  x"18",  x"00",  x"00",  x"3c",  x"3c", -- 02A0
         x"3e",  x"3f",  x"1f",  x"0c",  x"00",  x"00",  x"00",  x"00", -- 02A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"70", -- 02C8
         x"78",  x"7c",  x"3e",  x"3e",  x"3e",  x"1e",  x"00",  x"07", -- 02D0
         x"0f",  x"1f",  x"3e",  x"3e",  x"3e",  x"3c",  x"1e",  x"1e", -- 02D8
         x"3e",  x"3e",  x"3c",  x"18",  x"00",  x"00",  x"3c",  x"3c", -- 02E0
         x"3e",  x"3f",  x"1f",  x"0c",  x"00",  x"00",  x"00",  x"00", -- 02E8
         x"00",  x"00",  x"00",  x"1e",  x"1e",  x"0a",  x"00",  x"00", -- 02F0
         x"00",  x"00",  x"00",  x"3c",  x"3c",  x"28",  x"00",  x"00", -- 02F8
         x"10",  x"38",  x"18",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0300
         x"04",  x"0e",  x"0c",  x"00",  x"00",  x"00",  x"00",  x"50", -- 0308
         x"18",  x"5c",  x"30",  x"3f",  x"1e",  x"1b",  x"00",  x"05", -- 0310
         x"0c",  x"1d",  x"06",  x"7e",  x"3c",  x"6c",  x"00",  x"11", -- 0318
         x"10",  x"7d",  x"38",  x"08",  x"00",  x"00",  x"00",  x"44", -- 0320
         x"04",  x"5f",  x"0e",  x"08",  x"00",  x"00",  x"00",  x"00", -- 0328
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0330
         x"00",  x"06",  x"14",  x"18",  x"00",  x"00",  x"00",  x"00", -- 0338
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0340
         x"00",  x"00",  x"00",  x"01",  x"03",  x"07",  x"00",  x"00", -- 0348
         x"00",  x"00",  x"00",  x"00",  x"ff",  x"e0",  x"00",  x"00", -- 0350
         x"00",  x"00",  x"00",  x"00",  x"80",  x"c0",  x"07",  x"07", -- 0358
         x"00",  x"00",  x"00",  x"0f",  x"0f",  x"0f",  x"c0",  x"80", -- 0360
         x"01",  x"03",  x"3f",  x"ff",  x"ff",  x"ff",  x"c0",  x"e0", -- 0368
         x"e0",  x"f0",  x"f0",  x"f0",  x"f0",  x"f0",  x"07",  x"07", -- 0370
         x"04",  x"01",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff", -- 0378
         x"ff",  x"c3",  x"c3",  x"00",  x"00",  x"00",  x"e0",  x"e0", -- 0380
         x"c0",  x"80",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0388
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0390
         x"00",  x"60",  x"28",  x"18",  x"00",  x"00",  x"00",  x"00", -- 0398
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03A0
         x"00",  x"00",  x"00",  x"00",  x"01",  x"03",  x"00",  x"00", -- 03A8
         x"00",  x"00",  x"00",  x"00",  x"ff",  x"07",  x"00",  x"00", -- 03B0
         x"00",  x"00",  x"00",  x"80",  x"c0",  x"e0",  x"03",  x"07", -- 03B8
         x"07",  x"0f",  x"0f",  x"0f",  x"0f",  x"0f",  x"03",  x"01", -- 03C0
         x"80",  x"c0",  x"fc",  x"ff",  x"ff",  x"ff",  x"e0",  x"e0", -- 03C8
         x"00",  x"00",  x"00",  x"f0",  x"f0",  x"f0",  x"07",  x"07", -- 03D0
         x"03",  x"01",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff", -- 03D8
         x"ff",  x"c3",  x"c3",  x"00",  x"00",  x"00",  x"e0",  x"e0", -- 03E0
         x"20",  x"80",  x"5c",  x"01",  x"ff",  x"ff",  x"ff",  x"ff", -- 03E8
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 03F0
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
