library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_5800 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_5800;

architecture rtl of rom1_5800 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"06",  x"04",  x"3a",  x"35",  x"0d",  x"be",  x"28",  x"10", -- 0000
         x"1a",  x"77",  x"13",  x"23",  x"10",  x"f4",  x"af",  x"b9", -- 0008
         x"20",  x"0a",  x"01",  x"3c",  x"00",  x"09",  x"18",  x"e8", -- 0010
         x"d1",  x"c3",  x"86",  x"56",  x"21",  x"4b",  x"0d",  x"35", -- 0018
         x"28",  x"0f",  x"3e",  x"04",  x"be",  x"30",  x"11",  x"cb", -- 0020
         x"46",  x"28",  x"0d",  x"dd",  x"2b",  x"dd",  x"2b",  x"18", -- 0028
         x"0b",  x"ed",  x"5f",  x"e6",  x"0e",  x"c6",  x"04",  x"77", -- 0030
         x"dd",  x"23",  x"dd",  x"23",  x"d1",  x"c1",  x"e1",  x"c9", -- 0038
         x"21",  x"3c",  x"0d",  x"af",  x"be",  x"28",  x"f1",  x"3e", -- 0040
         x"3e",  x"be",  x"30",  x"01",  x"77",  x"11",  x"c0",  x"ff", -- 0048
         x"e5",  x"21",  x"50",  x"5c",  x"cd",  x"d4",  x"01",  x"e1", -- 0050
         x"eb",  x"3a",  x"3c",  x"0d",  x"85",  x"6f",  x"c5",  x"06", -- 0058
         x"08",  x"36",  x"dc",  x"23",  x"36",  x"de",  x"c5",  x"06", -- 0060
         x"08",  x"cd",  x"c7",  x"01",  x"10",  x"fb",  x"c1",  x"eb", -- 0068
         x"35",  x"eb",  x"28",  x"19",  x"36",  x"20",  x"2b",  x"36", -- 0070
         x"de",  x"2b",  x"36",  x"fc",  x"c5",  x"06",  x"05",  x"cd", -- 0078
         x"c7",  x"01",  x"10",  x"fb",  x"c1",  x"10",  x"da",  x"c1", -- 0080
         x"cd",  x"21",  x"59",  x"18",  x"ab",  x"2b",  x"2b",  x"36", -- 0088
         x"20",  x"23",  x"18",  x"f3",  x"c5",  x"e5",  x"06",  x"04", -- 0090
         x"36",  x"20",  x"23",  x"10",  x"fb",  x"01",  x"3f",  x"00", -- 0098
         x"09",  x"06",  x"04",  x"36",  x"20",  x"2b",  x"10",  x"fb", -- 00A0
         x"e1",  x"c1",  x"c9",  x"06",  x"08",  x"3e",  x"20",  x"be", -- 00A8
         x"c0",  x"23",  x"10",  x"fb",  x"3a",  x"46",  x"0d",  x"47", -- 00B0
         x"ed",  x"5f",  x"a0",  x"c0",  x"3a",  x"32",  x"0d",  x"fe", -- 00B8
         x"0f",  x"c0",  x"eb",  x"21",  x"40",  x"5c",  x"1b",  x"01", -- 00C0
         x"08",  x"00",  x"ed",  x"b8",  x"c9",  x"e5",  x"c5",  x"21", -- 00C8
         x"84",  x"f9",  x"0e",  x"0c",  x"db",  x"83",  x"cb",  x"5f", -- 00D0
         x"28",  x"1d",  x"e6",  x"07",  x"c6",  x"05",  x"47",  x"32", -- 00D8
         x"49",  x"0d",  x"3e",  x"50",  x"32",  x"4a",  x"0d",  x"36", -- 00E0
         x"d4",  x"23",  x"23",  x"cd",  x"41",  x"59",  x"21",  x"42", -- 00E8
         x"5c",  x"cd",  x"d4",  x"01",  x"c1",  x"e1",  x"c9",  x"cb", -- 00F0
         x"67",  x"28",  x"df",  x"36",  x"ce",  x"3e",  x"f4",  x"32", -- 00F8
         x"49",  x"0d",  x"3e",  x"50",  x"32",  x"4a",  x"0d",  x"06", -- 0100
         x"0c",  x"18",  x"de",  x"e5",  x"c5",  x"21",  x"84",  x"f9", -- 0108
         x"06",  x"0e",  x"36",  x"20",  x"23",  x"10",  x"fb",  x"c1", -- 0110
         x"e1",  x"af",  x"32",  x"49",  x"0d",  x"32",  x"4a",  x"0d", -- 0118
         x"c9",  x"e5",  x"c5",  x"21",  x"2c",  x"f8",  x"22",  x"3f", -- 0120
         x"0c",  x"2a",  x"3c",  x"0d",  x"22",  x"3d",  x"0c",  x"cd", -- 0128
         x"70",  x"02",  x"21",  x"c0",  x"ff",  x"3a",  x"3c",  x"0d", -- 0130
         x"47",  x"0e",  x"40",  x"cd",  x"41",  x"59",  x"c1",  x"e1", -- 0138
         x"c9",  x"af",  x"b8",  x"79",  x"28",  x"06",  x"90",  x"36", -- 0140
         x"d2",  x"23",  x"10",  x"fb",  x"47",  x"b7",  x"c8",  x"36", -- 0148
         x"20",  x"23",  x"10",  x"fb",  x"c9",  x"c5",  x"e5",  x"06", -- 0150
         x"20",  x"21",  x"02",  x"0d",  x"36",  x"00",  x"23",  x"10", -- 0158
         x"fb",  x"e1",  x"c1",  x"c9",  x"e5",  x"e5",  x"dd",  x"e1", -- 0160
         x"21",  x"00",  x"00",  x"22",  x"22",  x"0d",  x"7a",  x"01", -- 0168
         x"06",  x"00",  x"21",  x"39",  x"5b",  x"ed",  x"b1",  x"20", -- 0170
         x"2e",  x"7b",  x"e6",  x"70",  x"28",  x"12",  x"fe",  x"20", -- 0178
         x"28",  x"1a",  x"fe",  x"30",  x"28",  x"10",  x"fe",  x"50", -- 0180
         x"20",  x"1d",  x"3e",  x"10",  x"0e",  x"06",  x"18",  x"10", -- 0188
         x"3e",  x"58",  x"0e",  x"60",  x"18",  x"0a",  x"3e",  x"40", -- 0190
         x"0e",  x"60",  x"18",  x"04",  x"3e",  x"48",  x"0e",  x"06", -- 0198
         x"32",  x"22",  x"0d",  x"79",  x"32",  x"23",  x"0d",  x"21", -- 01A0
         x"02",  x"0d",  x"06",  x"08",  x"dd",  x"7e",  x"f8",  x"4e", -- 01A8
         x"cb",  x"3f",  x"cb",  x"19",  x"cb",  x"3f",  x"cb",  x"19", -- 01B0
         x"cb",  x"3f",  x"cb",  x"19",  x"cb",  x"3f",  x"cb",  x"19", -- 01B8
         x"71",  x"f5",  x"79",  x"17",  x"17",  x"17",  x"17",  x"e6", -- 01C0
         x"f0",  x"4f",  x"f1",  x"b1",  x"12",  x"d5",  x"4f",  x"3a", -- 01C8
         x"22",  x"0d",  x"83",  x"5f",  x"7a",  x"e6",  x"fe",  x"fe", -- 01D0
         x"f0",  x"79",  x"20",  x"04",  x"3a",  x"23",  x"0d",  x"b1", -- 01D8
         x"12",  x"d1",  x"23",  x"13",  x"dd",  x"23",  x"10",  x"c4", -- 01E0
         x"e1",  x"c9",  x"e5",  x"d5",  x"c5",  x"3e",  x"60",  x"21", -- 01E8
         x"60",  x"f0",  x"0e",  x"20",  x"11",  x"60",  x"00",  x"06", -- 01F0
         x"04",  x"c5",  x"41",  x"77",  x"23",  x"10",  x"fc",  x"19", -- 01F8
         x"c1",  x"10",  x"f6",  x"fe",  x"60",  x"28",  x"04",  x"c1", -- 0200
         x"d1",  x"e1",  x"c9",  x"21",  x"68",  x"f0",  x"0e",  x"10", -- 0208
         x"3e",  x"06",  x"11",  x"70",  x"00",  x"18",  x"e0",  x"00", -- 0210
         x"f8",  x"3f",  x"3d",  x"3d",  x"52",  x"45",  x"4b",  x"4f", -- 0218
         x"52",  x"44",  x"3a",  x"20",  x"30",  x"30",  x"20",  x"3d", -- 0220
         x"3d",  x"3d",  x"3d",  x"3d",  x"50",  x"55",  x"4e",  x"4b", -- 0228
         x"54",  x"45",  x"3a",  x"20",  x"30",  x"30",  x"20",  x"3d", -- 0230
         x"3d",  x"3d",  x"3d",  x"3d",  x"4d",  x"55",  x"4e",  x"49", -- 0238
         x"54",  x"49",  x"4f",  x"4e",  x"3a",  x"20",  x"30",  x"30", -- 0240
         x"20",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d", -- 0248
         x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d",  x"3d", -- 0250
         x"3d",  x"18",  x"f9",  x"0e",  x"4d",  x"55",  x"4c",  x"54", -- 0258
         x"49",  x"50",  x"4c",  x"49",  x"4b",  x"41",  x"54",  x"4f", -- 0260
         x"52",  x"3a",  x"0c",  x"fc",  x"1f",  x"4b",  x"45",  x"49", -- 0268
         x"4e",  x"45",  x"20",  x"4d",  x"55",  x"4e",  x"49",  x"54", -- 0270
         x"49",  x"4f",  x"4e",  x"20",  x"4d",  x"45",  x"48",  x"52", -- 0278
         x"20",  x"2d",  x"20",  x"53",  x"50",  x"49",  x"45",  x"4c", -- 0280
         x"45",  x"4e",  x"44",  x"45",  x"16",  x"fc",  x"0c",  x"4e", -- 0288
         x"45",  x"55",  x"45",  x"52",  x"20",  x"52",  x"45",  x"4b", -- 0290
         x"4f",  x"52",  x"44",  x"c7",  x"fc",  x"0a",  x"2d",  x"20", -- 0298
         x"20",  x"31",  x"20",  x"50",  x"55",  x"4e",  x"4b",  x"54", -- 02A0
         x"87",  x"fd",  x"0b",  x"2d",  x"20",  x"20",  x"32",  x"20", -- 02A8
         x"50",  x"55",  x"4e",  x"4b",  x"54",  x"45",  x"47",  x"fe", -- 02B0
         x"0b",  x"2d",  x"20",  x"20",  x"33",  x"20",  x"50",  x"55", -- 02B8
         x"4e",  x"4b",  x"54",  x"45",  x"d7",  x"fb",  x"11",  x"54", -- 02C0
         x"52",  x"45",  x"46",  x"46",  x"45",  x"52",  x"42",  x"45", -- 02C8
         x"57",  x"45",  x"52",  x"54",  x"55",  x"4e",  x"47",  x"3a", -- 02D0
         x"a5",  x"fc",  x"1a",  x"2d",  x"20",  x"20",  x"4d",  x"55", -- 02D8
         x"4e",  x"49",  x"54",  x"49",  x"4f",  x"4e",  x"20",  x"4a", -- 02E0
         x"45",  x"20",  x"4e",  x"41",  x"43",  x"48",  x"20",  x"49", -- 02E8
         x"4e",  x"48",  x"41",  x"4c",  x"54",  x"68",  x"fd",  x"15", -- 02F0
         x"5a",  x"49",  x"45",  x"4c",  x"46",  x"45",  x"4c",  x"44", -- 02F8
         x"45",  x"52",  x"20",  x"2d",  x"20",  x"45",  x"52",  x"48", -- 0300
         x"4f",  x"45",  x"48",  x"45",  x"4e",  x"a8",  x"fd",  x"12", -- 0308
         x"44",  x"45",  x"53",  x"20",  x"4d",  x"55",  x"4c",  x"54", -- 0310
         x"49",  x"50",  x"4c",  x"49",  x"4b",  x"41",  x"54",  x"4f", -- 0318
         x"52",  x"53",  x"e8",  x"fd",  x"14",  x"44",  x"45",  x"52", -- 0320
         x"20",  x"4a",  x"45",  x"57",  x"45",  x"49",  x"4c",  x"49", -- 0328
         x"47",  x"45",  x"4e",  x"20",  x"52",  x"45",  x"49",  x"48", -- 0330
         x"45",  x"ed",  x"ec",  x"f1",  x"f0",  x"f5",  x"f4",  x"06", -- 0338
         x"08",  x"09",  x"0b",  x"06",  x"08",  x"07",  x"09",  x"80", -- 0340
         x"a0",  x"00",  x"80",  x"a0",  x"b0",  x"80",  x"b0",  x"80", -- 0348
         x"80",  x"b0",  x"80",  x"b0",  x"b0",  x"80",  x"81",  x"81", -- 0350
         x"b1",  x"00",  x"00",  x"81",  x"81",  x"91",  x"b1",  x"b1", -- 0358
         x"81",  x"b1",  x"81",  x"b1",  x"81",  x"a0",  x"80",  x"b0", -- 0360
         x"00",  x"80",  x"00",  x"b0",  x"00",  x"00",  x"80",  x"80", -- 0368
         x"b0",  x"80",  x"00",  x"80",  x"8f",  x"01",  x"3f",  x"e9", -- 0370
         x"87",  x"01",  x"10",  x"00",  x"87",  x"01",  x"10",  x"e9", -- 0378
         x"87",  x"01",  x"10",  x"c4",  x"87",  x"01",  x"3f",  x"93", -- 0380
         x"87",  x"01",  x"10",  x"9c",  x"87",  x"01",  x"10",  x"93", -- 0388
         x"87",  x"01",  x"10",  x"83",  x"87",  x"01",  x"10",  x"93", -- 0390
         x"87",  x"01",  x"10",  x"9c",  x"87",  x"01",  x"10",  x"93", -- 0398
         x"87",  x"01",  x"10",  x"e9",  x"87",  x"01",  x"10",  x"c4", -- 03A0
         x"87",  x"01",  x"3f",  x"9c",  x"20",  x"9c",  x"00",  x"00", -- 03A8
         x"30",  x"dc",  x"87",  x"01",  x"10",  x"e9",  x"87",  x"01", -- 03B0
         x"10",  x"dc",  x"87",  x"01",  x"10",  x"af",  x"87",  x"01", -- 03B8
         x"3f",  x"9c",  x"87",  x"01",  x"20",  x"a5",  x"87",  x"01", -- 03C0
         x"10",  x"9c",  x"87",  x"01",  x"10",  x"93",  x"87",  x"01", -- 03C8
         x"10",  x"9c",  x"87",  x"01",  x"10",  x"a5",  x"87",  x"01", -- 03D0
         x"10",  x"9c",  x"87",  x"01",  x"10",  x"dc",  x"87",  x"01", -- 03D8
         x"10",  x"9c",  x"87",  x"01",  x"3f",  x"e9",  x"20",  x"e9", -- 03E0
         x"00",  x"e6",  x"e8",  x"ea",  x"20",  x"ec",  x"ee",  x"f0", -- 03E8
         x"20",  x"dc",  x"de",  x"20",  x"20",  x"20",  x"e0",  x"e2", -- 03F0
         x"e4",  x"fc",  x"de",  x"f2",  x"f4",  x"20",  x"e0",  x"e2"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
