library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_zre_0800 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom_zre_0800;

architecture rtl of rom_zre_0800 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"18",  x"2a",  x"18",  x"09",  x"f5",  x"3e",  x"03",  x"d3", -- 0000
         x"82",  x"f1",  x"c3",  x"62",  x"02",  x"f5",  x"e5",  x"2a", -- 0008
         x"80",  x"0f",  x"2b",  x"22",  x"80",  x"0f",  x"7c",  x"b5", -- 0010
         x"28",  x"05",  x"e1",  x"f1",  x"fb",  x"ed",  x"4d",  x"3e", -- 0018
         x"03",  x"d3",  x"82",  x"31",  x"ff",  x"0f",  x"21",  x"f1", -- 0020
         x"00",  x"e5",  x"18",  x"f0",  x"cd",  x"b7",  x"02",  x"21", -- 0028
         x"06",  x"f4",  x"11",  x"06",  x"ec",  x"06",  x"0c",  x"3e", -- 0030
         x"ff",  x"77",  x"12",  x"23",  x"13",  x"10",  x"fa",  x"21", -- 0038
         x"18",  x"ec",  x"11",  x"18",  x"f0",  x"06",  x"08",  x"77", -- 0040
         x"12",  x"23",  x"13",  x"10",  x"fa",  x"67",  x"6f",  x"22", -- 0048
         x"20",  x"ec",  x"21",  x"00",  x"00",  x"22",  x"20",  x"f4", -- 0050
         x"06",  x"20",  x"11",  x"3f",  x"00",  x"21",  x"00",  x"f8", -- 0058
         x"e5",  x"36",  x"83",  x"19",  x"36",  x"83",  x"23",  x"10", -- 0060
         x"f8",  x"e1",  x"cd",  x"d4",  x"09",  x"21",  x"40",  x"fa", -- 0068
         x"cd",  x"d4",  x"09",  x"21",  x"c0",  x"ff",  x"cd",  x"d4", -- 0070
         x"09",  x"21",  x"0b",  x"0a",  x"11",  x"96",  x"f8",  x"0e", -- 0078
         x"17",  x"ed",  x"b0",  x"11",  x"0d",  x"f9",  x"0e",  x"29", -- 0080
         x"ed",  x"b0",  x"1e",  x"4d",  x"0e",  x"28",  x"ed",  x"b0", -- 0088
         x"1e",  x"8d",  x"0e",  x"28",  x"ed",  x"b0",  x"1e",  x"d6", -- 0090
         x"0e",  x"16",  x"ed",  x"b0",  x"11",  x"d5",  x"fa",  x"0e", -- 0098
         x"17",  x"ed",  x"b0",  x"21",  x"15",  x"fb",  x"06",  x"17", -- 00A0
         x"36",  x"84",  x"23",  x"10",  x"fb",  x"11",  x"99",  x"fb", -- 00A8
         x"fd",  x"21",  x"50",  x"0f",  x"dd",  x"21",  x"ff",  x"01", -- 00B0
         x"d5",  x"16",  x"00",  x"dd",  x"5c",  x"21",  x"c7",  x"0a", -- 00B8
         x"19",  x"66",  x"fd",  x"74",  x"00",  x"6a",  x"5a",  x"42", -- 00C0
         x"4e",  x"eb",  x"09",  x"eb",  x"2c",  x"20",  x"f9",  x"dd", -- 00C8
         x"7c",  x"21",  x"be",  x"0a",  x"01",  x"13",  x"00",  x"09", -- 00D0
         x"3d",  x"20",  x"fc",  x"e5",  x"7e",  x"23",  x"66",  x"6f", -- 00D8
         x"97",  x"ed",  x"52",  x"e1",  x"28",  x"08",  x"2b",  x"7e", -- 00E0
         x"a7",  x"20",  x"e6",  x"d1",  x"18",  x"27",  x"d1",  x"dd", -- 00E8
         x"2c",  x"23",  x"23",  x"7e",  x"fd",  x"77",  x"01",  x"fd", -- 00F0
         x"23",  x"fd",  x"23",  x"23",  x"d5",  x"01",  x"0f",  x"00", -- 00F8
         x"ed",  x"b0",  x"d1",  x"3a",  x"02",  x"0c",  x"dd",  x"bd", -- 0100
         x"20",  x"06",  x"eb",  x"cd",  x"a2",  x"09",  x"e5",  x"eb", -- 0108
         x"21",  x"80",  x"00",  x"19",  x"eb",  x"dd",  x"24",  x"dd", -- 0110
         x"7c",  x"fe",  x"09",  x"20",  x"9b",  x"e1",  x"cd",  x"8f", -- 0118
         x"01",  x"f6",  x"e0",  x"fe",  x"ff",  x"28",  x"f7",  x"cb", -- 0120
         x"5f",  x"28",  x"43",  x"cb",  x"67",  x"28",  x"66",  x"cb", -- 0128
         x"47",  x"20",  x"eb",  x"21",  x"17",  x"fb",  x"11",  x"80", -- 0130
         x"00",  x"3e",  x"ff",  x"19",  x"3c",  x"cb",  x"7e",  x"28", -- 0138
         x"fa",  x"32",  x"02",  x"0c",  x"3c",  x"21",  x"4f",  x"0f", -- 0140
         x"23",  x"23",  x"3d",  x"20",  x"fb",  x"5e",  x"2b",  x"66", -- 0148
         x"6f",  x"3a",  x"03",  x"0c",  x"fe",  x"55",  x"28",  x"14", -- 0150
         x"e5",  x"65",  x"55",  x"06",  x"28",  x"19",  x"10",  x"fd", -- 0158
         x"22",  x"80",  x"0f",  x"e1",  x"3e",  x"b5",  x"d3",  x"82", -- 0160
         x"3e",  x"f4",  x"d3",  x"82",  x"f1",  x"e9",  x"e5",  x"11", -- 0168
         x"80",  x"ff",  x"19",  x"7e",  x"fe",  x"01",  x"e1",  x"fa", -- 0170
         x"1e",  x"09",  x"d5",  x"cd",  x"a0",  x"09",  x"d1",  x"19", -- 0178
         x"cd",  x"a2",  x"09",  x"11",  x"9b",  x"09",  x"eb",  x"cd", -- 0180
         x"e0",  x"01",  x"eb",  x"11",  x"00",  x"7f",  x"1b",  x"7a", -- 0188
         x"b3",  x"20",  x"fb",  x"18",  x"89",  x"e5",  x"11",  x"80", -- 0190
         x"00",  x"18",  x"d7",  x"01",  x"d8",  x"01",  x"00",  x"00", -- 0198
         x"97",  x"11",  x"3e",  x"81",  x"e5",  x"2b",  x"06",  x"03", -- 01A0
         x"2b",  x"77",  x"10",  x"fc",  x"a7",  x"28",  x"01",  x"3d", -- 01A8
         x"11",  x"41",  x"00",  x"ed",  x"52",  x"06",  x"17",  x"23", -- 01B0
         x"77",  x"10",  x"fc",  x"a7",  x"28",  x"01",  x"3c",  x"19", -- 01B8
         x"06",  x"03",  x"2b",  x"77",  x"10",  x"fc",  x"a7",  x"28", -- 01C0
         x"01",  x"3c",  x"23",  x"19",  x"06",  x"17",  x"77",  x"2b", -- 01C8
         x"10",  x"fc",  x"e1",  x"c9",  x"06",  x"40",  x"36",  x"83", -- 01D0
         x"23",  x"10",  x"fb",  x"c9",  x"00",  x"00",  x"00",  x"00", -- 01D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0200
         x"00",  x"00",  x"00",  x"57",  x"41",  x"45",  x"48",  x"4c", -- 0208
         x"45",  x"4e",  x"20",  x"53",  x"49",  x"45",  x"20",  x"49", -- 0210
         x"48",  x"52",  x"20",  x"53",  x"50",  x"49",  x"45",  x"4c", -- 0218
         x"20",  x"21",  x"44",  x"75",  x"72",  x"63",  x"68",  x"20", -- 0220
         x"41",  x"75",  x"66",  x"2d",  x"20",  x"75",  x"6e",  x"64", -- 0228
         x"20",  x"41",  x"62",  x"62",  x"65",  x"77",  x"65",  x"67", -- 0230
         x"75",  x"6e",  x"67",  x"20",  x"64",  x"65",  x"73",  x"20", -- 0238
         x"53",  x"70",  x"69",  x"65",  x"6c",  x"68",  x"65",  x"62", -- 0240
         x"65",  x"6c",  x"73",  x"77",  x"69",  x"72",  x"64",  x"20", -- 0248
         x"65",  x"69",  x"6e",  x"20",  x"53",  x"70",  x"69",  x"65", -- 0250
         x"6c",  x"20",  x"61",  x"75",  x"73",  x"67",  x"65",  x"73", -- 0258
         x"75",  x"63",  x"68",  x"74",  x"2e",  x"20",  x"4e",  x"61", -- 0260
         x"63",  x"68",  x"20",  x"44",  x"72",  x"75",  x"65",  x"63", -- 0268
         x"6b",  x"65",  x"6e",  x"64",  x"65",  x"73",  x"20",  x"53", -- 0270
         x"70",  x"69",  x"65",  x"6c",  x"6b",  x"6e",  x"6f",  x"70", -- 0278
         x"66",  x"65",  x"73",  x"20",  x"65",  x"72",  x"73",  x"63", -- 0280
         x"68",  x"65",  x"69",  x"6e",  x"74",  x"20",  x"64",  x"61", -- 0288
         x"73",  x"20",  x"76",  x"6f",  x"6e",  x"20",  x"49",  x"68", -- 0290
         x"6e",  x"65",  x"6e",  x"20",  x"20",  x"20",  x"67",  x"65", -- 0298
         x"77",  x"61",  x"65",  x"68",  x"6c",  x"74",  x"65",  x"20", -- 02A0
         x"53",  x"70",  x"69",  x"65",  x"6c",  x"2e",  x"20",  x"20", -- 02A8
         x"20",  x"53",  x"20",  x"50",  x"20",  x"49",  x"20",  x"45", -- 02B0
         x"20",  x"4c",  x"20",  x"41",  x"20",  x"55",  x"20",  x"53", -- 02B8
         x"20",  x"57",  x"20",  x"41",  x"20",  x"48",  x"20",  x"4c", -- 02C0
         x"1c",  x"28",  x"10",  x"40",  x"50",  x"60",  x"74",  x"80", -- 02C8
         x"00",  x"5c",  x"52",  x"14",  x"20",  x"20",  x"48",  x"49", -- 02D0
         x"52",  x"53",  x"43",  x"48",  x"4a",  x"41",  x"47",  x"44", -- 02D8
         x"20",  x"20",  x"20",  x"00",  x"d6",  x"55",  x"10",  x"20", -- 02E0
         x"48",  x"41",  x"53",  x"45",  x"20",  x"55",  x"4e",  x"44", -- 02E8
         x"20",  x"57",  x"4f",  x"4c",  x"46",  x"20",  x"0b",  x"b6", -- 02F0
         x"5a",  x"20",  x"20",  x"41",  x"42",  x"46",  x"41",  x"48", -- 02F8
         x"52",  x"54",  x"53",  x"4c",  x"41",  x"55",  x"46",  x"20", -- 0300
         x"20",  x"0a",  x"5c",  x"65",  x"0c",  x"53",  x"43",  x"48", -- 0308
         x"4d",  x"45",  x"54",  x"54",  x"45",  x"52",  x"4c",  x"49", -- 0310
         x"4e",  x"47",  x"45",  x"20",  x"00",  x"f1",  x"4e",  x"0f", -- 0318
         x"20",  x"20",  x"53",  x"43",  x"48",  x"49",  x"45",  x"53", -- 0320
         x"53",  x"42",  x"55",  x"44",  x"45",  x"20",  x"20",  x"0c", -- 0328
         x"0b",  x"54",  x"10",  x"20",  x"20",  x"41",  x"55",  x"54", -- 0330
         x"4f",  x"52",  x"45",  x"4e",  x"4e",  x"45",  x"4e",  x"20", -- 0338
         x"20",  x"20",  x"00",  x"f7",  x"5d",  x"1c",  x"20",  x"20", -- 0340
         x"20",  x"4d",  x"45",  x"52",  x"4b",  x"53",  x"50",  x"49", -- 0348
         x"45",  x"4c",  x"20",  x"20",  x"20",  x"09",  x"44",  x"37", -- 0350
         x"20",  x"57",  x"41",  x"53",  x"53",  x"45",  x"52",  x"52", -- 0358
         x"4f",  x"48",  x"52",  x"42",  x"52",  x"55",  x"43",  x"48", -- 0360
         x"00",  x"31",  x"5a",  x"20",  x"20",  x"44",  x"45",  x"52", -- 0368
         x"20",  x"47",  x"41",  x"45",  x"52",  x"54",  x"4e",  x"45", -- 0370
         x"52",  x"20",  x"20",  x"00",  x"bb",  x"29",  x"20",  x"49", -- 0378
         x"4d",  x"20",  x"47",  x"45",  x"57",  x"41",  x"45",  x"43", -- 0380
         x"48",  x"53",  x"48",  x"41",  x"55",  x"53",  x"00",  x"bd", -- 0388
         x"50",  x"1f",  x"48",  x"41",  x"47",  x"45",  x"4c",  x"4e", -- 0390
         x"44",  x"45",  x"20",  x"57",  x"4f",  x"4c",  x"4b",  x"45", -- 0398
         x"4e",  x"00",  x"71",  x"56",  x"20",  x"20",  x"20",  x"44", -- 03A0
         x"45",  x"52",  x"20",  x"54",  x"41",  x"55",  x"43",  x"48", -- 03A8
         x"45",  x"52",  x"20",  x"20",  x"00",  x"00",  x"00",  x"00", -- 03B0
         x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20", -- 03B8
         x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"00", -- 03C0
         x"00",  x"00",  x"00",  x"20",  x"20",  x"20",  x"20",  x"20", -- 03C8
         x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20", -- 03D0
         x"20",  x"20",  x"00",  x"00",  x"00",  x"00",  x"20",  x"20", -- 03D8
         x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20", -- 03E0
         x"20",  x"20",  x"20",  x"20",  x"20",  x"00",  x"00",  x"00", -- 03E8
         x"00",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20", -- 03F0
         x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20",  x"20"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
