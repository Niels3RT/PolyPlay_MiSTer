library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_6800 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_6800;

architecture rtl of rom1_6800 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"48",  x"57",  x"49",  x"4e",  x"44",  x"49",  x"47",  x"4b", -- 0000
         x"45",  x"49",  x"54",  x"20",  x"2b",  x"20",  x"46",  x"41", -- 0008
         x"48",  x"52",  x"54",  x"52",  x"49",  x"43",  x"48",  x"54", -- 0010
         x"55",  x"4e",  x"47",  x"29",  x"c9",  x"fb",  x"2e",  x"2d", -- 0018
         x"20",  x"47",  x"45",  x"47",  x"45",  x"4e",  x"53",  x"50", -- 0020
         x"49",  x"45",  x"4c",  x"45",  x"52",  x"20",  x"2d",  x"20", -- 0028
         x"52",  x"45",  x"43",  x"48",  x"4e",  x"45",  x"52",  x"47", -- 0030
         x"45",  x"53",  x"54",  x"45",  x"55",  x"45",  x"52",  x"54", -- 0038
         x"20",  x"28",  x"4c",  x"45",  x"52",  x"4e",  x"46",  x"41", -- 0040
         x"45",  x"48",  x"49",  x"47",  x"29",  x"04",  x"fd",  x"37", -- 0048
         x"45",  x"53",  x"20",  x"57",  x"45",  x"52",  x"44",  x"45", -- 0050
         x"4e",  x"20",  x"32",  x"20",  x"52",  x"45",  x"4e",  x"4e", -- 0058
         x"45",  x"4e",  x"20",  x"4d",  x"49",  x"54",  x"20",  x"4a", -- 0060
         x"45",  x"20",  x"34",  x"20",  x"52",  x"55",  x"4e",  x"44", -- 0068
         x"45",  x"4e",  x"20",  x"47",  x"45",  x"46",  x"41",  x"48", -- 0070
         x"52",  x"45",  x"4e",  x"2e",  x"20",  x"44",  x"45",  x"52", -- 0078
         x"20",  x"53",  x"49",  x"45",  x"47",  x"45",  x"52",  x"84", -- 0080
         x"fd",  x"39",  x"45",  x"52",  x"48",  x"41",  x"45",  x"4c", -- 0088
         x"54",  x"20",  x"46",  x"55",  x"45",  x"52",  x"20",  x"44", -- 0090
         x"41",  x"53",  x"20",  x"47",  x"45",  x"57",  x"4f",  x"4e", -- 0098
         x"4e",  x"45",  x"4e",  x"45",  x"20",  x"52",  x"45",  x"4e", -- 00A0
         x"4e",  x"45",  x"4e",  x"20",  x"44",  x"49",  x"45",  x"20", -- 00A8
         x"44",  x"4f",  x"50",  x"50",  x"45",  x"4c",  x"54",  x"45", -- 00B0
         x"20",  x"50",  x"55",  x"4e",  x"4b",  x"54",  x"5a",  x"41", -- 00B8
         x"48",  x"4c",  x"2e",  x"20",  x"93",  x"82",  x"01",  x"20", -- 00C0
         x"80",  x"bf",  x"01",  x"20",  x"93",  x"82",  x"01",  x"20", -- 00C8
         x"80",  x"ff",  x"01",  x"00",  x"3f",  x"ff",  x"00",  x"01", -- 00D0
         x"80",  x"00",  x"8f",  x"01",  x"48",  x"12",  x"82",  x"01", -- 00D8
         x"08",  x"e9",  x"82",  x"01",  x"08",  x"c4",  x"82",  x"01", -- 00E0
         x"20",  x"93",  x"00",  x"8f",  x"01",  x"08",  x"93",  x"82", -- 00E8
         x"01",  x"08",  x"c4",  x"82",  x"01",  x"08",  x"e9",  x"82", -- 00F0
         x"01",  x"60",  x"12",  x"00",  x"bf",  x"00",  x"08",  x"80", -- 00F8
         x"02",  x"60",  x"00",  x"8e",  x"00",  x"9c",  x"00",  x"80", -- 0100
         x"00",  x"aa",  x"00",  x"8e",  x"38",  x"9c",  x"38",  x"80", -- 0108
         x"38",  x"aa",  x"38",  x"01",  x"00",  x"c1",  x"ff",  x"c0", -- 0110
         x"ff",  x"bf",  x"ff",  x"ff",  x"ff",  x"3f",  x"00",  x"40", -- 0118
         x"00",  x"41",  x"00",  x"0b",  x"00",  x"09",  x"0e",  x"09", -- 0120
         x"02",  x"1f",  x"00",  x"02",  x"0e",  x"0a",  x"0c",  x"02", -- 0128
         x"0a",  x"17",  x"08",  x"17",  x"00",  x"02",  x"0e",  x"0a", -- 0130
         x"0c",  x"02",  x"0a",  x"1f",  x"08",  x"09",  x"06",  x"09", -- 0138
         x"0a",  x"0a",  x"08",  x"02",  x"06",  x"18",  x"04",  x"02", -- 0140
         x"02",  x"00",  x"16",  x"08",  x"07",  x"0a",  x"07",  x"0e", -- 0148
         x"15",  x"00",  x"00",  x"06",  x"0e",  x"05",  x"0a",  x"01", -- 0150
         x"08",  x"0a",  x"04",  x"00",  x"04",  x"0e",  x"00",  x"04", -- 0158
         x"02",  x"00",  x"04",  x"02",  x"00",  x"04",  x"0e",  x"00", -- 0160
         x"04",  x"0a",  x"00",  x"04",  x"06",  x"00",  x"04",  x"06", -- 0168
         x"00",  x"04",  x"0a",  x"00",  x"0b",  x"0e",  x"02",  x"00", -- 0170
         x"0a",  x"02",  x"00",  x"05",  x"0e",  x"04",  x"0c",  x"04", -- 0178
         x"0a",  x"00",  x"05",  x"0a",  x"04",  x"0c",  x"04",  x"0e", -- 0180
         x"00",  x"05",  x"0e",  x"04",  x"0c",  x"04",  x"0a",  x"00", -- 0188
         x"0b",  x"06",  x"02",  x"08",  x"0a",  x"0a",  x"00",  x"07", -- 0190
         x"08",  x"02",  x"0a",  x"10",  x"0c",  x"02",  x"0e",  x"05", -- 0198
         x"00",  x"00",  x"03",  x"0e",  x"00",  x"03",  x"06",  x"00", -- 01A0
         x"03",  x"02",  x"00",  x"03",  x"0a",  x"00",  x"04",  x"0e", -- 01A8
         x"02",  x"0a",  x"02",  x"0c",  x"03",  x"02",  x"04",  x"0c", -- 01B0
         x"01",  x"00",  x"02",  x"04",  x"01",  x"0e",  x"05",  x"00", -- 01B8
         x"00",  x"04",  x"02",  x"02",  x"06",  x"02",  x"04",  x"03", -- 01C0
         x"0e",  x"04",  x"04",  x"01",  x"00",  x"02",  x"0c",  x"01", -- 01C8
         x"02",  x"05",  x"00",  x"00",  x"f6",  x"f8",  x"a2",  x"69", -- 01D0
         x"e2",  x"ff",  x"a5",  x"69",  x"f6",  x"ff",  x"a8",  x"69", -- 01D8
         x"e2",  x"f8",  x"ab",  x"69",  x"c0",  x"fc",  x"ae",  x"69", -- 01E0
         x"c0",  x"fb",  x"c1",  x"69",  x"0c",  x"0e",  x"0a",  x"1a", -- 01E8
         x"12",  x"16",  x"14",  x"1c",  x"10",  x"c4",  x"87",  x"01", -- 01F0
         x"18",  x"c4",  x"8f",  x"01",  x"10",  x"c4",  x"87",  x"01", -- 01F8
         x"10",  x"d0",  x"87",  x"01",  x"10",  x"c4",  x"87",  x"01", -- 0200
         x"10",  x"af",  x"87",  x"01",  x"10",  x"c4",  x"87",  x"01", -- 0208
         x"10",  x"75",  x"87",  x"01",  x"18",  x"75",  x"8f",  x"01", -- 0210
         x"10",  x"93",  x"87",  x"01",  x"30",  x"c4",  x"ff",  x"01", -- 0218
         x"00",  x"00",  x"00",  x"11",  x"00",  x"00",  x"00",  x"00", -- 0220
         x"00",  x"00",  x"00",  x"3c",  x"00",  x"00",  x"00",  x"00", -- 0228
         x"00",  x"39",  x"7f",  x"ff",  x"00",  x"00",  x"00",  x"00", -- 0230
         x"00",  x"c0",  x"e0",  x"f3",  x"00",  x"00",  x"00",  x"00", -- 0238
         x"00",  x"00",  x"00",  x"c0",  x"3c",  x"3c",  x"3c",  x"3c", -- 0240
         x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"f9",  x"e0", -- 0248
         x"e0",  x"c0",  x"c0",  x"e0",  x"f3",  x"f3",  x"f3",  x"73", -- 0250
         x"70",  x"30",  x"30",  x"70",  x"c0",  x"c0",  x"c0",  x"c0", -- 0258
         x"00",  x"00",  x"00",  x"00",  x"3c",  x"3c",  x"3c",  x"3c", -- 0260
         x"3c",  x"00",  x"00",  x"00",  x"e0",  x"f9",  x"ff",  x"ff", -- 0268
         x"ff",  x"7f",  x"39",  x"00",  x"73",  x"f3",  x"f3",  x"f3", -- 0270
         x"f3",  x"e0",  x"c0",  x"00",  x"c0",  x"c0",  x"c0",  x"c0", -- 0278
         x"c0",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"f9",  x"e0", -- 0280
         x"e0",  x"c0",  x"c0",  x"e0",  x"f3",  x"f3",  x"f3",  x"73", -- 0288
         x"70",  x"30",  x"30",  x"70",  x"00",  x"00",  x"00",  x"00", -- 0290
         x"00",  x"0f",  x"0f",  x"0f",  x"00",  x"00",  x"00",  x"00", -- 0298
         x"00",  x"e0",  x"e0",  x"e0",  x"00",  x"00",  x"00",  x"00", -- 02A0
         x"00",  x"7f",  x"7f",  x"7f",  x"08",  x"00",  x"0d",  x"00", -- 02A8
         x"00",  x"1f",  x"3f",  x"7f",  x"3f",  x"3f",  x"7f",  x"00", -- 02B0
         x"00",  x"ff",  x"f9",  x"c0",  x"00",  x"00",  x"c0",  x"00", -- 02B8
         x"00",  x"ff",  x"ff",  x"3f",  x"0f",  x"0f",  x"3f",  x"00", -- 02C0
         x"00",  x"80",  x"c0",  x"e0",  x"c0",  x"c0",  x"e0",  x"3f", -- 02C8
         x"1f",  x"00",  x"00",  x"0f",  x"0f",  x"0f",  x"00",  x"f9", -- 02D0
         x"ff",  x"00",  x"00",  x"e0",  x"e0",  x"e0",  x"00",  x"ff", -- 02D8
         x"ff",  x"00",  x"00",  x"7f",  x"7f",  x"7f",  x"00",  x"c0", -- 02E0
         x"80",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02E8
         x"00",  x"ff",  x"f9",  x"c0",  x"00",  x"00",  x"c0",  x"00", -- 02F0
         x"00",  x"ff",  x"ff",  x"3f",  x"0f",  x"0f",  x"3f",  x"00", -- 02F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"01",  x"00",  x"00", -- 0300
         x"00",  x"00",  x"18",  x"7c",  x"fe",  x"f8",  x"f3",  x"00", -- 0308
         x"00",  x"00",  x"00",  x"00",  x"00",  x"f8",  x"fe",  x"08", -- 0310
         x"00",  x"0a",  x"00",  x"10",  x"78",  x"fc",  x"f8",  x"e7", -- 0318
         x"47",  x"1f",  x"27",  x"0f",  x"3f",  x"78",  x"f8",  x"f0", -- 0320
         x"81",  x"c3",  x"ff",  x"ff",  x"ff",  x"3f",  x"3f",  x"3e", -- 0328
         x"fc",  x"f1",  x"00",  x"80",  x"80",  x"80",  x"80",  x"40", -- 0330
         x"f0",  x"f8",  x"1f",  x"1f",  x"1f",  x"0f",  x"07",  x"03", -- 0338
         x"00",  x"00",  x"c3",  x"ff",  x"ff",  x"fc",  x"f8",  x"f3", -- 0340
         x"07",  x"0f",  x"e7",  x"c3",  x"00",  x"40",  x"e0",  x"f0", -- 0348
         x"e0",  x"c0",  x"f0",  x"c0",  x"80",  x"00",  x"00",  x"00", -- 0350
         x"00",  x"00",  x"27",  x"0f",  x"3f",  x"78",  x"f8",  x"f0", -- 0358
         x"81",  x"c3",  x"ff",  x"ff",  x"ff",  x"3f",  x"3f",  x"3e", -- 0360
         x"fc",  x"f1",  x"08",  x"00",  x"1b",  x"00",  x"00",  x"00", -- 0368
         x"00",  x"00",  x"00",  x"1f",  x"7f",  x"00",  x"00",  x"00", -- 0370
         x"18",  x"3e",  x"7f",  x"1f",  x"0f",  x"00",  x"00",  x"00", -- 0378
         x"00",  x"00",  x"00",  x"80",  x"00",  x"00",  x"01",  x"01", -- 0380
         x"01",  x"01",  x"04",  x"0f",  x"1f",  x"ff",  x"ff",  x"ff", -- 0388
         x"fc",  x"fc",  x"ec",  x"3f",  x"0e",  x"e4",  x"f0",  x"fc", -- 0390
         x"16",  x"03",  x"07",  x"01",  x"03",  x"00",  x"08",  x"1e", -- 0398
         x"3f",  x"1f",  x"e7",  x"e2",  x"f8",  x"0f",  x"03",  x"01", -- 03A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"e7",  x"c3",  x"00", -- 03A8
         x"02",  x"07",  x"0f",  x"07",  x"03",  x"c3",  x"ff",  x"ff", -- 03B0
         x"3f",  x"1f",  x"cf",  x"e0",  x"f0",  x"f8",  x"f8",  x"f8", -- 03B8
         x"f0",  x"e0",  x"c0",  x"00",  x"00",  x"ff",  x"ff",  x"ff", -- 03C0
         x"fc",  x"fc",  x"ec",  x"3f",  x"0e",  x"e4",  x"f0",  x"fc", -- 03C8
         x"16",  x"03",  x"07",  x"01",  x"03",  x"00",  x"00",  x"00", -- 03D0
         x"3c",  x"3c",  x"3c",  x"3c",  x"3c",  x"00",  x"39",  x"7f", -- 03D8
         x"ff",  x"ff",  x"ff",  x"f9",  x"e0",  x"00",  x"c0",  x"e0", -- 03E0
         x"f3",  x"f3",  x"f3",  x"f3",  x"73",  x"00",  x"00",  x"00", -- 03E8
         x"c0",  x"c0",  x"c0",  x"c0",  x"c0",  x"00",  x"00",  x"00", -- 03F0
         x"00",  x"3c",  x"3c",  x"3c",  x"3c",  x"e0",  x"c0",  x"c0"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
