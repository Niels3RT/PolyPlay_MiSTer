library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_5400 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_5400;

architecture rtl of rom1_5400 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"da",  x"54",  x"5d",  x"13",  x"01",  x"3f",  x"02",  x"ed", -- 0000
         x"b0",  x"2a",  x"18",  x"0c",  x"ed",  x"5b",  x"0c",  x"0c", -- 0008
         x"b7",  x"ed",  x"52",  x"38",  x"14",  x"cd",  x"0b",  x"57", -- 0010
         x"8c",  x"5a",  x"2a",  x"18",  x"0c",  x"22",  x"0c",  x"0c", -- 0018
         x"21",  x"74",  x"5b",  x"cd",  x"e0",  x"01",  x"c3",  x"f1", -- 0020
         x"00",  x"cd",  x"0b",  x"57",  x"6a",  x"5a",  x"18",  x"f0", -- 0028
         x"c5",  x"d5",  x"3a",  x"00",  x"0d",  x"3d",  x"28",  x"19", -- 0030
         x"3e",  x"7f",  x"11",  x"40",  x"00",  x"06",  x"3c",  x"be", -- 0038
         x"30",  x"01",  x"34",  x"19",  x"be",  x"30",  x"01",  x"34", -- 0040
         x"37",  x"ed",  x"52",  x"10",  x"f2",  x"b7",  x"d1",  x"c1", -- 0048
         x"c9",  x"e5",  x"f5",  x"3a",  x"32",  x"0d",  x"83",  x"5f", -- 0050
         x"30",  x"01",  x"14",  x"ed",  x"a8",  x"c5",  x"01",  x"41", -- 0058
         x"00",  x"09",  x"c1",  x"ed",  x"a8",  x"f1",  x"e1",  x"06", -- 0060
         x"3b",  x"11",  x"3f",  x"00",  x"2b",  x"7e",  x"e6",  x"fe", -- 0068
         x"23",  x"77",  x"19",  x"7e",  x"e6",  x"fe",  x"23",  x"77", -- 0070
         x"37",  x"ed",  x"52",  x"2b",  x"2b",  x"10",  x"ee",  x"23", -- 0078
         x"37",  x"d1",  x"c1",  x"c9",  x"c5",  x"d5",  x"3a",  x"00", -- 0080
         x"0d",  x"3d",  x"28",  x"1f",  x"3e",  x"7f",  x"11",  x"40", -- 0088
         x"00",  x"06",  x"3c",  x"be",  x"30",  x"01",  x"35",  x"19", -- 0090
         x"be",  x"30",  x"01",  x"35",  x"b7",  x"23",  x"ed",  x"52", -- 0098
         x"10",  x"f1",  x"b7",  x"d1",  x"c1",  x"f5",  x"cd",  x"6f", -- 00A0
         x"57",  x"f1",  x"c9",  x"e5",  x"f5",  x"3a",  x"32",  x"0d", -- 00A8
         x"83",  x"5f",  x"30",  x"01",  x"14",  x"ed",  x"a8",  x"c5", -- 00B0
         x"01",  x"41",  x"00",  x"09",  x"c1",  x"ed",  x"a8",  x"f1", -- 00B8
         x"e1",  x"06",  x"3b",  x"11",  x"41",  x"00",  x"23",  x"7e", -- 00C0
         x"fe",  x"7f",  x"38",  x"02",  x"f6",  x"01",  x"2b",  x"77", -- 00C8
         x"19",  x"7e",  x"fe",  x"7f",  x"38",  x"02",  x"f6",  x"01", -- 00D0
         x"2b",  x"77",  x"b7",  x"ed",  x"52",  x"23",  x"23",  x"23", -- 00D8
         x"10",  x"e5",  x"2b",  x"37",  x"d1",  x"c1",  x"f5",  x"cd", -- 00E0
         x"6f",  x"57",  x"f1",  x"c9",  x"eb",  x"23",  x"3a",  x"33", -- 00E8
         x"0d",  x"85",  x"6f",  x"30",  x"01",  x"24",  x"ed",  x"a8", -- 00F0
         x"eb",  x"c5",  x"01",  x"41",  x"00",  x"09",  x"c1",  x"eb", -- 00F8
         x"ed",  x"a0",  x"c9",  x"3a",  x"32",  x"0d",  x"83",  x"5f", -- 0100
         x"30",  x"01",  x"14",  x"1a",  x"e6",  x"fe",  x"77",  x"c5", -- 0108
         x"01",  x"40",  x"00",  x"09",  x"c1",  x"1b",  x"1a",  x"e6", -- 0110
         x"fe",  x"77",  x"c9",  x"06",  x"0f",  x"1a",  x"b7",  x"28", -- 0118
         x"03",  x"cd",  x"79",  x"55",  x"cd",  x"c7",  x"01",  x"13", -- 0120
         x"23",  x"23",  x"23",  x"23",  x"10",  x"ef",  x"c9",  x"e5", -- 0128
         x"2a",  x"39",  x"0d",  x"3e",  x"77",  x"bd",  x"38",  x"11", -- 0130
         x"3a",  x"35",  x"0d",  x"cb",  x"47",  x"20",  x"0e",  x"36", -- 0138
         x"c3",  x"23",  x"36",  x"c5",  x"3e",  x"c1",  x"32",  x"35", -- 0140
         x"0d",  x"3e",  x"ff",  x"e1",  x"c9",  x"36",  x"20",  x"23", -- 0148
         x"22",  x"39",  x"0d",  x"36",  x"c2",  x"23",  x"36",  x"c4", -- 0150
         x"3e",  x"c0",  x"32",  x"35",  x"0d",  x"18",  x"ea",  x"e5", -- 0158
         x"2a",  x"39",  x"0d",  x"3e",  x"42",  x"bd",  x"28",  x"e1", -- 0160
         x"3a",  x"35",  x"0d",  x"cb",  x"47",  x"20",  x"e4",  x"23", -- 0168
         x"36",  x"20",  x"2b",  x"2b",  x"22",  x"39",  x"0d",  x"18", -- 0170
         x"c6",  x"d5",  x"f5",  x"e5",  x"c5",  x"11",  x"3d",  x"00", -- 0178
         x"01",  x"01",  x"03",  x"77",  x"c6",  x"02",  x"23",  x"10", -- 0180
         x"fa",  x"0d",  x"20",  x"05",  x"06",  x"03",  x"19",  x"18", -- 0188
         x"f2",  x"c1",  x"e1",  x"f1",  x"d1",  x"c9",  x"e5",  x"c5", -- 0190
         x"fd",  x"cb",  x"00",  x"46",  x"28",  x"0b",  x"db",  x"84", -- 0198
         x"1f",  x"1f",  x"d4",  x"2f",  x"55",  x"1f",  x"d4",  x"5f", -- 01A0
         x"55",  x"cd",  x"c7",  x"01",  x"21",  x"34",  x"0d",  x"35", -- 01A8
         x"28",  x"52",  x"2a",  x"37",  x"0d",  x"3a",  x"3b",  x"0d", -- 01B0
         x"77",  x"01",  x"c0",  x"ff",  x"09",  x"7e",  x"32",  x"3b", -- 01B8
         x"0d",  x"fe",  x"c6",  x"d2",  x"6b",  x"56",  x"fe",  x"10", -- 01C0
         x"ca",  x"90",  x"56",  x"fe",  x"80",  x"38",  x"2b",  x"e5", -- 01C8
         x"01",  x"04",  x"00",  x"e6",  x"0f",  x"21",  x"35",  x"0d", -- 01D0
         x"cb",  x"46",  x"28",  x"05",  x"21",  x"43",  x"5b",  x"18", -- 01D8
         x"03",  x"21",  x"3f",  x"5b",  x"ed",  x"b1",  x"e1",  x"28", -- 01E0
         x"24",  x"cb",  x"47",  x"28",  x"0d",  x"47",  x"3a",  x"3b", -- 01E8
         x"0d",  x"cb",  x"18",  x"e6",  x"f0",  x"f6",  x"0c",  x"b0", -- 01F0
         x"18",  x"03",  x"3a",  x"36",  x"0d",  x"77",  x"22",  x"37", -- 01F8
         x"0d",  x"c1",  x"e1",  x"c9",  x"34",  x"2a",  x"37",  x"0d", -- 0200
         x"36",  x"20",  x"c1",  x"e1",  x"c9",  x"06",  x"03",  x"c5", -- 0208
         x"d6",  x"06",  x"cb",  x"2f",  x"28",  x"04",  x"2b",  x"3d", -- 0210
         x"20",  x"fc",  x"36",  x"20",  x"23",  x"10",  x"fb",  x"2b", -- 0218
         x"01",  x"c0",  x"ff",  x"09",  x"c1",  x"7e",  x"36",  x"20", -- 0220
         x"2b",  x"10",  x"fb",  x"0e",  x"02",  x"fe",  x"90",  x"38", -- 0228
         x"07",  x"0d",  x"fe",  x"b0",  x"38",  x"02",  x"0e",  x"03", -- 0230
         x"21",  x"3f",  x"0d",  x"3a",  x"34",  x"0d",  x"d6",  x"10", -- 0238
         x"28",  x"03",  x"30",  x"02",  x"23",  x"23",  x"7e",  x"e5", -- 0240
         x"2a",  x"18",  x"0c",  x"85",  x"6f",  x"30",  x"01",  x"24", -- 0248
         x"22",  x"18",  x"0c",  x"22",  x"3d",  x"0c",  x"e1",  x"0d", -- 0250
         x"20",  x"ec",  x"21",  x"1a",  x"f8",  x"22",  x"3f",  x"0c", -- 0258
         x"cd",  x"70",  x"02",  x"21",  x"49",  x"5c",  x"cd",  x"d4", -- 0260
         x"01",  x"18",  x"25",  x"fe",  x"d0",  x"28",  x"68",  x"fe", -- 0268
         x"c8",  x"28",  x"87",  x"fe",  x"da",  x"28",  x"27",  x"fe", -- 0270
         x"d6",  x"28",  x"33",  x"fe",  x"d8",  x"28",  x"3f",  x"3a", -- 0278
         x"34",  x"0d",  x"fe",  x"14",  x"38",  x"0a",  x"2a",  x"47", -- 0280
         x"0d",  x"cd",  x"94",  x"58",  x"dd",  x"21",  x"37",  x"5c", -- 0288
         x"3e",  x"01",  x"32",  x"34",  x"0d",  x"21",  x"7e",  x"f9", -- 0290
         x"22",  x"37",  x"0d",  x"c1",  x"e1",  x"c9",  x"21",  x"3f", -- 0298
         x"0d",  x"34",  x"7e",  x"21",  x"78",  x"f9",  x"cd",  x"2a", -- 02A0
         x"57",  x"21",  x"ff",  x"fc",  x"18",  x"1e",  x"21",  x"40", -- 02A8
         x"0d",  x"34",  x"7e",  x"21",  x"72",  x"f9",  x"cd",  x"2a", -- 02B0
         x"57",  x"21",  x"3f",  x"fc",  x"18",  x"0e",  x"21",  x"41", -- 02B8
         x"0d",  x"34",  x"7e",  x"21",  x"6c",  x"f9",  x"cd",  x"2a", -- 02C0
         x"57",  x"21",  x"7f",  x"fb",  x"cd",  x"2a",  x"57",  x"21", -- 02C8
         x"5f",  x"5c",  x"cd",  x"d4",  x"01",  x"18",  x"b9",  x"3a", -- 02D0
         x"49",  x"0d",  x"fe",  x"00",  x"28",  x"b2",  x"f5",  x"fa", -- 02D8
         x"ea",  x"56",  x"21",  x"5f",  x"5c",  x"cd",  x"d4",  x"01", -- 02E0
         x"18",  x"06",  x"21",  x"50",  x"5c",  x"cd",  x"e0",  x"01", -- 02E8
         x"f1",  x"21",  x"3c",  x"0d",  x"86",  x"77",  x"f2",  x"03", -- 02F0
         x"57",  x"36",  x"00",  x"cd",  x"21",  x"59",  x"cd",  x"0b", -- 02F8
         x"59",  x"18",  x"8d",  x"fe",  x"41",  x"38",  x"f4",  x"36", -- 0300
         x"40",  x"18",  x"f0",  x"e1",  x"5e",  x"23",  x"56",  x"23", -- 0308
         x"e5",  x"d5",  x"e1",  x"5e",  x"23",  x"56",  x"23",  x"4e", -- 0310
         x"06",  x"00",  x"23",  x"ed",  x"b0",  x"c9",  x"c5",  x"06", -- 0318
         x"08",  x"7e",  x"b1",  x"12",  x"23",  x"13",  x"10",  x"f9", -- 0320
         x"c1",  x"c9",  x"e5",  x"c5",  x"f5",  x"f5",  x"01",  x"c0", -- 0328
         x"ff",  x"09",  x"06",  x"00",  x"04",  x"d6",  x"0a",  x"30", -- 0330
         x"fb",  x"f1",  x"c6",  x"06",  x"10",  x"fc",  x"d6",  x"06", -- 0338
         x"47",  x"e6",  x"0f",  x"c6",  x"30",  x"77",  x"78",  x"1f", -- 0340
         x"1f",  x"1f",  x"1f",  x"2b",  x"e6",  x"0f",  x"28",  x"03", -- 0348
         x"c6",  x"30",  x"77",  x"f1",  x"c1",  x"e1",  x"c9",  x"e5", -- 0350
         x"21",  x"42",  x"0d",  x"35",  x"20",  x"0f",  x"36",  x"08", -- 0358
         x"23",  x"ed",  x"5f",  x"e6",  x"03",  x"28",  x"04",  x"36", -- 0360
         x"c8",  x"18",  x"02",  x"36",  x"c6",  x"e1",  x"c9",  x"e5", -- 0368
         x"c5",  x"21",  x"d7",  x"f9",  x"cd",  x"57",  x"57",  x"cb", -- 0370
         x"46",  x"20",  x"47",  x"3a",  x"43",  x"0d",  x"77",  x"7e", -- 0378
         x"06",  x"28",  x"23",  x"be",  x"28",  x"19",  x"7e",  x"cb", -- 0380
         x"47",  x"20",  x"07",  x"f6",  x"01",  x"77",  x"e6",  x"fe", -- 0388
         x"18",  x"0d",  x"f5",  x"2f",  x"e6",  x"0f",  x"4f",  x"f1", -- 0390
         x"e6",  x"f0",  x"b1",  x"77",  x"23",  x"7e",  x"2b",  x"10", -- 0398
         x"e1",  x"01",  x"40",  x"00",  x"7e",  x"09",  x"06",  x"28", -- 03A0
         x"cb",  x"47",  x"20",  x"01",  x"77",  x"7e",  x"2b",  x"be", -- 03A8
         x"28",  x"0e",  x"cb",  x"46",  x"28",  x"05",  x"7e",  x"e6", -- 03B0
         x"fe",  x"18",  x"01",  x"3c",  x"77",  x"2b",  x"7e",  x"23", -- 03B8
         x"10",  x"ec",  x"c1",  x"e1",  x"c9",  x"dd",  x"cb",  x"01", -- 03C0
         x"76",  x"c0",  x"e5",  x"c5",  x"d5",  x"3a",  x"59",  x"0c", -- 03C8
         x"b7",  x"20",  x"06",  x"21",  x"66",  x"5c",  x"cd",  x"d4", -- 03D0
         x"01",  x"dd",  x"5e",  x"00",  x"16",  x"00",  x"cb",  x"7b", -- 03D8
         x"28",  x"01",  x"15",  x"2a",  x"47",  x"0d",  x"cd",  x"94", -- 03E0
         x"58",  x"dd",  x"cb",  x"01",  x"7e",  x"20",  x"51",  x"19", -- 03E8
         x"22",  x"47",  x"0d",  x"11",  x"e9",  x"5b",  x"dd",  x"7e", -- 03F0
         x"01",  x"83",  x"5f",  x"30",  x"01",  x"14",  x"0e",  x"00"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
