library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom1_8000 is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end rom1_8000;

architecture rtl of rom1_8000 is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"cd",  x"8f",  x"8b",  x"c3",  x"c9",  x"83",  x"07",  x"0f", -- 0000
         x"1a",  x"1f",  x"1f",  x"0d",  x"07",  x"00",  x"00",  x"00", -- 0008
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"06",  x"0c", -- 0010
         x"0c",  x"0c",  x"18",  x"18",  x"30",  x"00",  x"c0",  x"c0", -- 0018
         x"60",  x"60",  x"c0",  x"80",  x"80",  x"00",  x"0c",  x"0c", -- 0020
         x"18",  x"18",  x"0c",  x"06",  x"06",  x"00",  x"80",  x"c0", -- 0028
         x"c0",  x"c0",  x"60",  x"60",  x"30",  x"00",  x"06",  x"02", -- 0030
         x"02",  x"02",  x"03",  x"00",  x"00",  x"00",  x"0c",  x"08", -- 0038
         x"08",  x"08",  x"f8",  x"00",  x"00",  x"00",  x"06",  x"02", -- 0040
         x"02",  x"02",  x"03",  x"00",  x"00",  x"00",  x"0c",  x"08", -- 0048
         x"08",  x"08",  x"f8",  x"00",  x"00",  x"00",  x"06",  x"02", -- 0050
         x"02",  x"02",  x"03",  x"00",  x"00",  x"00",  x"0c",  x"08", -- 0058
         x"08",  x"08",  x"f8",  x"00",  x"00",  x"00",  x"c0",  x"c0", -- 0060
         x"80",  x"80",  x"80",  x"80",  x"80",  x"00",  x"31",  x"1b", -- 0068
         x"0e",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0070
         x"0f",  x"9f",  x"df",  x"4f",  x"9f",  x"c6",  x"00",  x"00", -- 0078
         x"00",  x"80",  x"80",  x"80",  x"00",  x"00",  x"00",  x"88", -- 0080
         x"c8",  x"c8",  x"cc",  x"c8",  x"84",  x"04",  x"00",  x"02", -- 0088
         x"02",  x"02",  x"06",  x"04",  x"04",  x"04",  x"00",  x"88", -- 0090
         x"c8",  x"c8",  x"cc",  x"c8",  x"84",  x"04",  x"00",  x"02", -- 0098
         x"02",  x"02",  x"06",  x"04",  x"04",  x"04",  x"00",  x"88", -- 00A0
         x"c8",  x"c8",  x"cc",  x"c8",  x"84",  x"04",  x"00",  x"02", -- 00A8
         x"02",  x"02",  x"06",  x"04",  x"04",  x"04",  x"00",  x"88", -- 00B0
         x"c8",  x"c8",  x"cc",  x"c8",  x"84",  x"04",  x"00",  x"02", -- 00B8
         x"02",  x"02",  x"06",  x"04",  x"04",  x"04",  x"00",  x"88", -- 00C0
         x"c8",  x"c8",  x"cc",  x"c8",  x"84",  x"04",  x"00",  x"02", -- 00C8
         x"02",  x"02",  x"06",  x"04",  x"04",  x"04",  x"00",  x"00", -- 00D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 00D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"81",  x"81", -- 00E0
         x"01",  x"01",  x"01",  x"01",  x"81",  x"81",  x"81",  x"81", -- 00E8
         x"81",  x"81",  x"81",  x"81",  x"81",  x"81",  x"00",  x"0c", -- 00F0
         x"06",  x"03",  x"01",  x"80",  x"c0",  x"60",  x"18",  x"3c", -- 00F8
         x"3c",  x"38",  x"18",  x"00",  x"00",  x"00",  x"00",  x"0f", -- 0100
         x"1a",  x"1f",  x"18",  x"0f",  x"07",  x"1f",  x"3f",  x"3f", -- 0108
         x"3f",  x"3f",  x"3f",  x"3f",  x"3f",  x"1f",  x"00",  x"00", -- 0110
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0118
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0120
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0128
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"e0",  x"e0", -- 0130
         x"f8",  x"fc",  x"ec",  x"e0",  x"e0",  x"c0",  x"00",  x"00", -- 0138
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"e0",  x"e0", -- 0140
         x"f8",  x"fc",  x"ec",  x"e0",  x"e0",  x"c0",  x"00",  x"00", -- 0148
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"e0",  x"e0", -- 0150
         x"f8",  x"fc",  x"ec",  x"e0",  x"e0",  x"c0",  x"00",  x"00", -- 0158
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0160
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0168
         x"01",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0170
         x"0f",  x"1f",  x"1f",  x"1f",  x"0f",  x"06",  x"00",  x"00", -- 0178
         x"00",  x"80",  x"80",  x"80",  x"00",  x"00",  x"00",  x"00", -- 0180
         x"80",  x"c0",  x"c0",  x"c0",  x"80",  x"00",  x"00",  x"00", -- 0188
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0190
         x"80",  x"c0",  x"c0",  x"c0",  x"80",  x"00",  x"00",  x"00", -- 0198
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01A0
         x"80",  x"c0",  x"c0",  x"c0",  x"80",  x"00",  x"00",  x"00", -- 01A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01B0
         x"80",  x"c0",  x"c0",  x"c0",  x"80",  x"00",  x"00",  x"00", -- 01B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01C0
         x"80",  x"c0",  x"c0",  x"c0",  x"80",  x"00",  x"00",  x"00", -- 01C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"18",  x"3c", -- 01F8
         x"3c",  x"38",  x"18",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0200
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"aa",  x"aa", -- 0208
         x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"aa",  x"55", -- 0210
         x"aa",  x"55",  x"aa",  x"55",  x"aa",  x"55",  x"ff",  x"3f", -- 0218
         x"3f",  x"3f",  x"3f",  x"3f",  x"3f",  x"1f",  x"80",  x"c0", -- 0220
         x"c0",  x"c0",  x"c0",  x"c0",  x"c0",  x"80",  x"00",  x"00", -- 0228
         x"00",  x"00",  x"00",  x"00",  x"00",  x"ff",  x"00",  x"00", -- 0230
         x"00",  x"00",  x"00",  x"00",  x"ff",  x"ff",  x"00",  x"00", -- 0238
         x"00",  x"00",  x"00",  x"ff",  x"ff",  x"ff",  x"00",  x"00", -- 0240
         x"00",  x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"00", -- 0248
         x"00",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"00", -- 0250
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"ff", -- 0258
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff", -- 0260
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"00",  x"00", -- 0268
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0270
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"06",  x"0c", -- 0278
         x"0c",  x"0c",  x"18",  x"18",  x"30",  x"00",  x"c0",  x"c0", -- 0280
         x"60",  x"60",  x"c0",  x"80",  x"80",  x"00",  x"0c",  x"0c", -- 0288
         x"18",  x"18",  x"0c",  x"06",  x"06",  x"00",  x"80",  x"c0", -- 0290
         x"c0",  x"c0",  x"60",  x"60",  x"30",  x"00",  x"00",  x"00", -- 0298
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02A8
         x"01",  x"01",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02B0
         x"f0",  x"f0",  x"00",  x"00",  x"00",  x"00",  x"01",  x"01", -- 02B8
         x"01",  x"01",  x"00",  x"00",  x"00",  x"00",  x"f0",  x"f0", -- 02C0
         x"f0",  x"f0",  x"00",  x"00",  x"00",  x"00",  x"c0",  x"c0", -- 02C8
         x"80",  x"80",  x"80",  x"80",  x"80",  x"00",  x"00",  x"00", -- 02D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02F8
         x"00",  x"00",  x"00",  x"00",  x"03",  x"03",  x"00",  x"00", -- 0300
         x"00",  x"00",  x"00",  x"00",  x"f8",  x"f8",  x"00",  x"00", -- 0308
         x"00",  x"00",  x"03",  x"03",  x"03",  x"03",  x"00",  x"00", -- 0310
         x"00",  x"00",  x"f8",  x"f8",  x"f8",  x"f8",  x"00",  x"00", -- 0318
         x"07",  x"07",  x"03",  x"03",  x"03",  x"03",  x"00",  x"00", -- 0320
         x"fc",  x"fc",  x"f8",  x"f8",  x"f8",  x"f8",  x"1f",  x"17", -- 0328
         x"17",  x"07",  x"03",  x"03",  x"03",  x"03",  x"fe",  x"fc", -- 0330
         x"fc",  x"fc",  x"f8",  x"f8",  x"f8",  x"f8",  x"07",  x"0f", -- 0338
         x"3f",  x"7f",  x"ff",  x"ff",  x"ff",  x"ff",  x"0c",  x"3f", -- 0340
         x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"ff",  x"7e",  x"7e", -- 0348
         x"fe",  x"fe",  x"fe",  x"fe",  x"7e",  x"7e",  x"7e",  x"7e", -- 0350
         x"7e",  x"7e",  x"7e",  x"7e",  x"7e",  x"7e",  x"00",  x"00", -- 0358
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"18",  x"3c", -- 0360
         x"3c",  x"38",  x"18",  x"00",  x"00",  x"00",  x"10",  x"af", -- 0368
         x"82",  x"01",  x"10",  x"af",  x"82",  x"01",  x"10",  x"9c", -- 0370
         x"82",  x"01",  x"10",  x"9c",  x"82",  x"01",  x"20",  x"af", -- 0378
         x"82",  x"01",  x"00",  x"00",  x"10",  x"af",  x"82",  x"01", -- 0380
         x"10",  x"af",  x"82",  x"01",  x"10",  x"9c",  x"82",  x"01", -- 0388
         x"00",  x"08",  x"40",  x"08",  x"30",  x"08",  x"20",  x"00", -- 0390
         x"04",  x"28",  x"04",  x"38",  x"04",  x"48",  x"00",  x"10", -- 0398
         x"af",  x"82",  x"01",  x"10",  x"af",  x"82",  x"01",  x"20", -- 03A0
         x"83",  x"82",  x"01",  x"00",  x"08",  x"28",  x"08",  x"38", -- 03A8
         x"00",  x"08",  x"20",  x"08",  x"30",  x"08",  x"40",  x"08", -- 03B0
         x"50",  x"00",  x"18",  x"00",  x"82",  x"01",  x"08",  x"00", -- 03B8
         x"82",  x"01",  x"20",  x"c4",  x"82",  x"01",  x"20",  x"9c", -- 03C0
         x"00",  x"cd",  x"b7",  x"02",  x"21",  x"50",  x"00",  x"11", -- 03C8
         x"06",  x"80",  x"01",  x"00",  x"01",  x"cd",  x"c8",  x"02", -- 03D0
         x"21",  x"50",  x"00",  x"11",  x"06",  x"81",  x"01",  x"28", -- 03D8
         x"01",  x"cd",  x"ce",  x"02",  x"21",  x"48",  x"00",  x"11", -- 03E0
         x"2e",  x"82",  x"01",  x"40",  x"01",  x"cd",  x"d4",  x"02", -- 03E8
         x"cd",  x"53",  x"8b",  x"11",  x"d3",  x"f9",  x"21",  x"35", -- 03F0
         x"8c",  x"01",  x"1d",  x"00",  x"ed",  x"b0",  x"06",  x"06"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
